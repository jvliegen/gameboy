library IEEE;

use IEEE.STD_LOGIC_1164.ALL;

entity gameboy_v1 is
  port (
    reset : in STD_LOGIC;
    clock : in STD_LOGIC;

  );
end gameboy_v1;

architecture Behavioural of gameboy_v1 is

  signal reset_i, clock_i : STD_LOGIC;

begin
  
  -------------------------------------------------------------------------------
  -- (DE-)LOCALISING IN/OUTPUTS
  -------------------------------------------------------------------------------
  reset_i <= reset;
  clock_i <= clock;

  
  -------------------------------------------------------------------------------
  -- processor
  -------------------------------------------------------------------------------


  -------------------------------------------------------------------------------
  -- ROM
  -------------------------------------------------------------------------------


  -------------------------------------------------------------------------------
  -- RAM
  -------------------------------------------------------------------------------

end Behavioural;