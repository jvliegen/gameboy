library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library work;
use work.PKG_gameboy.ALL;

entity processor_tb is
end processor_tb;

architecture Behavioural of processor_tb is

  signal reset, clock : STD_LOGIC;

  signal bus_we : STD_LOGIC;
  signal bus_address : STD_LOGIC_VECTOR(15 downto 0);
  signal bus_data_in, bus_data_out : STD_LOGIC_VECTOR(7 downto 0);


  constant clock_period : time := 250 ns;

begin

  -------------------------------------------------------------------------------
  -- STIMULI
  -------------------------------------------------------------------------------
  PSTIM: process
  begin
    reset <= '1';
    wait for clock_period*2;

    reset <= '0';
    wait for clock_period*2;



    wait;
  end process;

  -------------------------------------------------------------------------------
  -- MEMORY MODEL
  -------------------------------------------------------------------------------
  PMUX: process(bus_address)
  begin
    case bus_address is
      when x"0040" => bus_data_in <= x"d9";
      when x"0048" => bus_data_in <= x"d9";
      when x"0050" => bus_data_in <= x"d9";
      when x"0058" => bus_data_in <= x"d9";
      when x"0060" => bus_data_in <= x"d9";
      when x"0061" => bus_data_in <= x"04";
      when x"0062" => bus_data_in <= x"0c";
      when x"0063" => bus_data_in <= x"18";
      when x"0064" => bus_data_in <= x"01";
      when x"0065" => bus_data_in <= x"22";
      when x"0066" => bus_data_in <= x"0d";
      when x"0067" => bus_data_in <= x"20";
      when x"0068" => bus_data_in <= x"fc";
      when x"0069" => bus_data_in <= x"05";
      when x"006a" => bus_data_in <= x"20";
      when x"006b" => bus_data_in <= x"f9";
      when x"006c" => bus_data_in <= x"c9";
      when x"006d" => bus_data_in <= x"04";
      when x"006e" => bus_data_in <= x"0c";
      when x"006f" => bus_data_in <= x"18";
      when x"0070" => bus_data_in <= x"03";
      when x"0071" => bus_data_in <= x"2a";
      when x"0072" => bus_data_in <= x"12";
      when x"0073" => bus_data_in <= x"13";
      when x"0074" => bus_data_in <= x"0d";
      when x"0075" => bus_data_in <= x"20";
      when x"0076" => bus_data_in <= x"fa";
      when x"0077" => bus_data_in <= x"05";
      when x"0078" => bus_data_in <= x"20";
      when x"0079" => bus_data_in <= x"f7";
      when x"007a" => bus_data_in <= x"c9";
      when x"007b" => bus_data_in <= x"04";
      when x"007c" => bus_data_in <= x"0c";
      when x"007d" => bus_data_in <= x"18";
      when x"007e" => bus_data_in <= x"05";
      when x"007f" => bus_data_in <= x"2a";
      when x"0080" => bus_data_in <= x"12";
      when x"0081" => bus_data_in <= x"13";
      when x"0082" => bus_data_in <= x"12";
      when x"0083" => bus_data_in <= x"13";
      when x"0084" => bus_data_in <= x"0d";
      when x"0085" => bus_data_in <= x"20";
      when x"0086" => bus_data_in <= x"f8";
      when x"0087" => bus_data_in <= x"05";
      when x"0088" => bus_data_in <= x"20";
      when x"0089" => bus_data_in <= x"f5";
      when x"008a" => bus_data_in <= x"c9";
      when x"008b" => bus_data_in <= x"04";
      when x"008c" => bus_data_in <= x"0c";
      when x"008d" => bus_data_in <= x"18";
      when x"008e" => bus_data_in <= x"0b";
      when x"008f" => bus_data_in <= x"f5";
      when x"0090" => bus_data_in <= x"f3";
      when x"0091" => bus_data_in <= x"f0";
      when x"0092" => bus_data_in <= x"41";
      when x"0093" => bus_data_in <= x"e6";
      when x"0094" => bus_data_in <= x"02";
      when x"0095" => bus_data_in <= x"20";
      when x"0096" => bus_data_in <= x"fa";
      when x"0097" => bus_data_in <= x"f1";
      when x"0098" => bus_data_in <= x"22";
      when x"0099" => bus_data_in <= x"fb";
      when x"009a" => bus_data_in <= x"0d";
      when x"009b" => bus_data_in <= x"20";
      when x"009c" => bus_data_in <= x"f2";
      when x"009d" => bus_data_in <= x"05";
      when x"009e" => bus_data_in <= x"20";
      when x"009f" => bus_data_in <= x"ef";
      when x"00a0" => bus_data_in <= x"c9";
      when x"00a1" => bus_data_in <= x"04";
      when x"00a2" => bus_data_in <= x"0c";
      when x"00a3" => bus_data_in <= x"18";
      when x"00a4" => bus_data_in <= x"0b";
      when x"00a5" => bus_data_in <= x"f3";
      when x"00a6" => bus_data_in <= x"f0";
      when x"00a7" => bus_data_in <= x"41";
      when x"00a8" => bus_data_in <= x"e6";
      when x"00a9" => bus_data_in <= x"02";
      when x"00aa" => bus_data_in <= x"20";
      when x"00ab" => bus_data_in <= x"fa";
      when x"00ac" => bus_data_in <= x"2a";
      when x"00ad" => bus_data_in <= x"12";
      when x"00ae" => bus_data_in <= x"fb";
      when x"00af" => bus_data_in <= x"13";
      when x"00b0" => bus_data_in <= x"0d";
      when x"00b1" => bus_data_in <= x"20";
      when x"00b2" => bus_data_in <= x"f2";
      when x"00b3" => bus_data_in <= x"05";
      when x"00b4" => bus_data_in <= x"20";
      when x"00b5" => bus_data_in <= x"ef";
      when x"00b6" => bus_data_in <= x"c9";
      when x"0101" => bus_data_in <= x"c3";
      when x"0102" => bus_data_in <= x"52";
      when x"0103" => bus_data_in <= x"09";
      when x"0104" => bus_data_in <= x"ce";
      when x"0105" => bus_data_in <= x"ed";
      when x"0106" => bus_data_in <= x"66";
      when x"0107" => bus_data_in <= x"66";
      when x"0108" => bus_data_in <= x"cc";
      when x"0109" => bus_data_in <= x"0d";
      when x"010b" => bus_data_in <= x"0b";
      when x"010c" => bus_data_in <= x"03";
      when x"010d" => bus_data_in <= x"73";
      when x"010f" => bus_data_in <= x"83";
      when x"0111" => bus_data_in <= x"0c";
      when x"0113" => bus_data_in <= x"0d";
      when x"0115" => bus_data_in <= x"08";
      when x"0116" => bus_data_in <= x"11";
      when x"0117" => bus_data_in <= x"1f";
      when x"0118" => bus_data_in <= x"88";
      when x"0119" => bus_data_in <= x"89";
      when x"011b" => bus_data_in <= x"0e";
      when x"011c" => bus_data_in <= x"dc";
      when x"011d" => bus_data_in <= x"cc";
      when x"011e" => bus_data_in <= x"6e";
      when x"011f" => bus_data_in <= x"e6";
      when x"0120" => bus_data_in <= x"dd";
      when x"0121" => bus_data_in <= x"dd";
      when x"0122" => bus_data_in <= x"d9";
      when x"0123" => bus_data_in <= x"99";
      when x"0124" => bus_data_in <= x"bb";
      when x"0125" => bus_data_in <= x"bb";
      when x"0126" => bus_data_in <= x"67";
      when x"0127" => bus_data_in <= x"63";
      when x"0128" => bus_data_in <= x"6e";
      when x"0129" => bus_data_in <= x"0e";
      when x"012a" => bus_data_in <= x"ec";
      when x"012b" => bus_data_in <= x"cc";
      when x"012c" => bus_data_in <= x"dd";
      when x"012d" => bus_data_in <= x"dc";
      when x"012e" => bus_data_in <= x"99";
      when x"012f" => bus_data_in <= x"9f";
      when x"0130" => bus_data_in <= x"bb";
      when x"0131" => bus_data_in <= x"b9";
      when x"0132" => bus_data_in <= x"33";
      when x"0133" => bus_data_in <= x"3e";
      when x"0134" => bus_data_in <= x"45";
      when x"0135" => bus_data_in <= x"58";
      when x"0136" => bus_data_in <= x"41";
      when x"0137" => bus_data_in <= x"4d";
      when x"0138" => bus_data_in <= x"50";
      when x"0139" => bus_data_in <= x"4c";
      when x"013a" => bus_data_in <= x"45";
      when x"014a" => bus_data_in <= x"01";
      when x"014b" => bus_data_in <= x"33";
      when x"014d" => bus_data_in <= x"a7";
      when x"014e" => bus_data_in <= x"f8";
      when x"014f" => bus_data_in <= x"5f";
      when x"0150" => bus_data_in <= x"7e";
      when x"0151" => bus_data_in <= x"42";
      when x"0152" => bus_data_in <= x"42";
      when x"0153" => bus_data_in <= x"42";
      when x"0154" => bus_data_in <= x"42";
      when x"0155" => bus_data_in <= x"42";
      when x"0156" => bus_data_in <= x"42";
      when x"0157" => bus_data_in <= x"7e";
      when x"0158" => bus_data_in <= x"7e";
      when x"0159" => bus_data_in <= x"81";
      when x"015a" => bus_data_in <= x"a5";
      when x"015b" => bus_data_in <= x"81";
      when x"015c" => bus_data_in <= x"bd";
      when x"015d" => bus_data_in <= x"99";
      when x"015e" => bus_data_in <= x"81";
      when x"015f" => bus_data_in <= x"7e";
      when x"0160" => bus_data_in <= x"7e";
      when x"0161" => bus_data_in <= x"ff";
      when x"0162" => bus_data_in <= x"db";
      when x"0163" => bus_data_in <= x"ff";
      when x"0164" => bus_data_in <= x"c3";
      when x"0165" => bus_data_in <= x"e7";
      when x"0166" => bus_data_in <= x"ff";
      when x"0167" => bus_data_in <= x"7e";
      when x"0168" => bus_data_in <= x"6c";
      when x"0169" => bus_data_in <= x"fe";
      when x"016a" => bus_data_in <= x"fe";
      when x"016b" => bus_data_in <= x"fe";
      when x"016c" => bus_data_in <= x"7c";
      when x"016d" => bus_data_in <= x"38";
      when x"016e" => bus_data_in <= x"10";
      when x"0170" => bus_data_in <= x"10";
      when x"0171" => bus_data_in <= x"38";
      when x"0172" => bus_data_in <= x"7c";
      when x"0173" => bus_data_in <= x"fe";
      when x"0174" => bus_data_in <= x"7c";
      when x"0175" => bus_data_in <= x"38";
      when x"0176" => bus_data_in <= x"10";
      when x"0178" => bus_data_in <= x"38";
      when x"0179" => bus_data_in <= x"7c";
      when x"017a" => bus_data_in <= x"38";
      when x"017b" => bus_data_in <= x"fe";
      when x"017c" => bus_data_in <= x"fe";
      when x"017d" => bus_data_in <= x"7c";
      when x"017e" => bus_data_in <= x"38";
      when x"017f" => bus_data_in <= x"7c";
      when x"0180" => bus_data_in <= x"10";
      when x"0181" => bus_data_in <= x"10";
      when x"0182" => bus_data_in <= x"38";
      when x"0183" => bus_data_in <= x"7c";
      when x"0184" => bus_data_in <= x"fe";
      when x"0185" => bus_data_in <= x"7c";
      when x"0186" => bus_data_in <= x"38";
      when x"0187" => bus_data_in <= x"7c";
      when x"018a" => bus_data_in <= x"18";
      when x"018b" => bus_data_in <= x"3c";
      when x"018c" => bus_data_in <= x"3c";
      when x"018d" => bus_data_in <= x"18";
      when x"0190" => bus_data_in <= x"ff";
      when x"0191" => bus_data_in <= x"ff";
      when x"0192" => bus_data_in <= x"e7";
      when x"0193" => bus_data_in <= x"c3";
      when x"0194" => bus_data_in <= x"c3";
      when x"0195" => bus_data_in <= x"e7";
      when x"0196" => bus_data_in <= x"ff";
      when x"0197" => bus_data_in <= x"ff";
      when x"0199" => bus_data_in <= x"3c";
      when x"019a" => bus_data_in <= x"66";
      when x"019b" => bus_data_in <= x"42";
      when x"019c" => bus_data_in <= x"42";
      when x"019d" => bus_data_in <= x"66";
      when x"019e" => bus_data_in <= x"3c";
      when x"01a0" => bus_data_in <= x"ff";
      when x"01a1" => bus_data_in <= x"c3";
      when x"01a2" => bus_data_in <= x"99";
      when x"01a3" => bus_data_in <= x"bd";
      when x"01a4" => bus_data_in <= x"bd";
      when x"01a5" => bus_data_in <= x"99";
      when x"01a6" => bus_data_in <= x"c3";
      when x"01a7" => bus_data_in <= x"ff";
      when x"01a8" => bus_data_in <= x"0f";
      when x"01a9" => bus_data_in <= x"07";
      when x"01aa" => bus_data_in <= x"0f";
      when x"01ab" => bus_data_in <= x"7d";
      when x"01ac" => bus_data_in <= x"cc";
      when x"01ad" => bus_data_in <= x"cc";
      when x"01ae" => bus_data_in <= x"cc";
      when x"01af" => bus_data_in <= x"78";
      when x"01b0" => bus_data_in <= x"3c";
      when x"01b1" => bus_data_in <= x"66";
      when x"01b2" => bus_data_in <= x"66";
      when x"01b3" => bus_data_in <= x"66";
      when x"01b4" => bus_data_in <= x"3c";
      when x"01b5" => bus_data_in <= x"18";
      when x"01b6" => bus_data_in <= x"7e";
      when x"01b7" => bus_data_in <= x"18";
      when x"01b8" => bus_data_in <= x"3f";
      when x"01b9" => bus_data_in <= x"33";
      when x"01ba" => bus_data_in <= x"3f";
      when x"01bb" => bus_data_in <= x"30";
      when x"01bc" => bus_data_in <= x"30";
      when x"01bd" => bus_data_in <= x"70";
      when x"01be" => bus_data_in <= x"f0";
      when x"01bf" => bus_data_in <= x"e0";
      when x"01c0" => bus_data_in <= x"7f";
      when x"01c1" => bus_data_in <= x"63";
      when x"01c2" => bus_data_in <= x"7f";
      when x"01c3" => bus_data_in <= x"63";
      when x"01c4" => bus_data_in <= x"63";
      when x"01c5" => bus_data_in <= x"67";
      when x"01c6" => bus_data_in <= x"e6";
      when x"01c7" => bus_data_in <= x"c0";
      when x"01c8" => bus_data_in <= x"99";
      when x"01c9" => bus_data_in <= x"5a";
      when x"01ca" => bus_data_in <= x"3c";
      when x"01cb" => bus_data_in <= x"e7";
      when x"01cc" => bus_data_in <= x"e7";
      when x"01cd" => bus_data_in <= x"3c";
      when x"01ce" => bus_data_in <= x"5a";
      when x"01cf" => bus_data_in <= x"99";
      when x"01d0" => bus_data_in <= x"80";
      when x"01d1" => bus_data_in <= x"e0";
      when x"01d2" => bus_data_in <= x"f8";
      when x"01d3" => bus_data_in <= x"fe";
      when x"01d4" => bus_data_in <= x"f8";
      when x"01d5" => bus_data_in <= x"e0";
      when x"01d6" => bus_data_in <= x"80";
      when x"01d8" => bus_data_in <= x"02";
      when x"01d9" => bus_data_in <= x"0e";
      when x"01da" => bus_data_in <= x"3e";
      when x"01db" => bus_data_in <= x"fe";
      when x"01dc" => bus_data_in <= x"3e";
      when x"01dd" => bus_data_in <= x"0e";
      when x"01de" => bus_data_in <= x"02";
      when x"01e0" => bus_data_in <= x"18";
      when x"01e1" => bus_data_in <= x"3c";
      when x"01e2" => bus_data_in <= x"7e";
      when x"01e3" => bus_data_in <= x"18";
      when x"01e4" => bus_data_in <= x"18";
      when x"01e5" => bus_data_in <= x"7e";
      when x"01e6" => bus_data_in <= x"3c";
      when x"01e7" => bus_data_in <= x"18";
      when x"01e8" => bus_data_in <= x"66";
      when x"01e9" => bus_data_in <= x"66";
      when x"01ea" => bus_data_in <= x"66";
      when x"01eb" => bus_data_in <= x"66";
      when x"01ec" => bus_data_in <= x"66";
      when x"01ee" => bus_data_in <= x"66";
      when x"01f0" => bus_data_in <= x"7f";
      when x"01f1" => bus_data_in <= x"db";
      when x"01f2" => bus_data_in <= x"db";
      when x"01f3" => bus_data_in <= x"7b";
      when x"01f4" => bus_data_in <= x"1b";
      when x"01f5" => bus_data_in <= x"1b";
      when x"01f6" => bus_data_in <= x"1b";
      when x"01f8" => bus_data_in <= x"3e";
      when x"01f9" => bus_data_in <= x"63";
      when x"01fa" => bus_data_in <= x"38";
      when x"01fb" => bus_data_in <= x"6c";
      when x"01fc" => bus_data_in <= x"6c";
      when x"01fd" => bus_data_in <= x"38";
      when x"01fe" => bus_data_in <= x"cc";
      when x"01ff" => bus_data_in <= x"78";
      when x"0204" => bus_data_in <= x"7e";
      when x"0205" => bus_data_in <= x"7e";
      when x"0206" => bus_data_in <= x"7e";
      when x"0208" => bus_data_in <= x"18";
      when x"0209" => bus_data_in <= x"3c";
      when x"020a" => bus_data_in <= x"7e";
      when x"020b" => bus_data_in <= x"18";
      when x"020c" => bus_data_in <= x"7e";
      when x"020d" => bus_data_in <= x"3c";
      when x"020e" => bus_data_in <= x"18";
      when x"020f" => bus_data_in <= x"ff";
      when x"0210" => bus_data_in <= x"18";
      when x"0211" => bus_data_in <= x"3c";
      when x"0212" => bus_data_in <= x"7e";
      when x"0213" => bus_data_in <= x"18";
      when x"0214" => bus_data_in <= x"18";
      when x"0215" => bus_data_in <= x"18";
      when x"0216" => bus_data_in <= x"18";
      when x"0218" => bus_data_in <= x"18";
      when x"0219" => bus_data_in <= x"18";
      when x"021a" => bus_data_in <= x"18";
      when x"021b" => bus_data_in <= x"18";
      when x"021c" => bus_data_in <= x"7e";
      when x"021d" => bus_data_in <= x"3c";
      when x"021e" => bus_data_in <= x"18";
      when x"0221" => bus_data_in <= x"18";
      when x"0222" => bus_data_in <= x"0c";
      when x"0223" => bus_data_in <= x"fe";
      when x"0224" => bus_data_in <= x"0c";
      when x"0225" => bus_data_in <= x"18";
      when x"0229" => bus_data_in <= x"30";
      when x"022a" => bus_data_in <= x"60";
      when x"022b" => bus_data_in <= x"fe";
      when x"022c" => bus_data_in <= x"60";
      when x"022d" => bus_data_in <= x"30";
      when x"0232" => bus_data_in <= x"c0";
      when x"0233" => bus_data_in <= x"c0";
      when x"0234" => bus_data_in <= x"c0";
      when x"0235" => bus_data_in <= x"fe";
      when x"0239" => bus_data_in <= x"24";
      when x"023a" => bus_data_in <= x"66";
      when x"023b" => bus_data_in <= x"ff";
      when x"023c" => bus_data_in <= x"66";
      when x"023d" => bus_data_in <= x"24";
      when x"0241" => bus_data_in <= x"18";
      when x"0242" => bus_data_in <= x"3c";
      when x"0243" => bus_data_in <= x"7e";
      when x"0244" => bus_data_in <= x"ff";
      when x"0245" => bus_data_in <= x"ff";
      when x"0249" => bus_data_in <= x"ff";
      when x"024a" => bus_data_in <= x"ff";
      when x"024b" => bus_data_in <= x"7e";
      when x"024c" => bus_data_in <= x"3c";
      when x"024d" => bus_data_in <= x"18";
      when x"0258" => bus_data_in <= x"30";
      when x"0259" => bus_data_in <= x"30";
      when x"025a" => bus_data_in <= x"30";
      when x"025b" => bus_data_in <= x"30";
      when x"025c" => bus_data_in <= x"30";
      when x"025e" => bus_data_in <= x"30";
      when x"0260" => bus_data_in <= x"6c";
      when x"0261" => bus_data_in <= x"6c";
      when x"0262" => bus_data_in <= x"6c";
      when x"0268" => bus_data_in <= x"6c";
      when x"0269" => bus_data_in <= x"6c";
      when x"026a" => bus_data_in <= x"fe";
      when x"026b" => bus_data_in <= x"6c";
      when x"026c" => bus_data_in <= x"fe";
      when x"026d" => bus_data_in <= x"6c";
      when x"026e" => bus_data_in <= x"6c";
      when x"0270" => bus_data_in <= x"30";
      when x"0271" => bus_data_in <= x"7c";
      when x"0272" => bus_data_in <= x"c0";
      when x"0273" => bus_data_in <= x"78";
      when x"0274" => bus_data_in <= x"0c";
      when x"0275" => bus_data_in <= x"f8";
      when x"0276" => bus_data_in <= x"30";
      when x"0279" => bus_data_in <= x"c6";
      when x"027a" => bus_data_in <= x"cc";
      when x"027b" => bus_data_in <= x"18";
      when x"027c" => bus_data_in <= x"30";
      when x"027d" => bus_data_in <= x"66";
      when x"027e" => bus_data_in <= x"c6";
      when x"0280" => bus_data_in <= x"38";
      when x"0281" => bus_data_in <= x"6c";
      when x"0282" => bus_data_in <= x"38";
      when x"0283" => bus_data_in <= x"76";
      when x"0284" => bus_data_in <= x"dc";
      when x"0285" => bus_data_in <= x"cc";
      when x"0286" => bus_data_in <= x"76";
      when x"0288" => bus_data_in <= x"60";
      when x"0289" => bus_data_in <= x"60";
      when x"028a" => bus_data_in <= x"c0";
      when x"0290" => bus_data_in <= x"18";
      when x"0291" => bus_data_in <= x"30";
      when x"0292" => bus_data_in <= x"60";
      when x"0293" => bus_data_in <= x"60";
      when x"0294" => bus_data_in <= x"60";
      when x"0295" => bus_data_in <= x"30";
      when x"0296" => bus_data_in <= x"18";
      when x"0298" => bus_data_in <= x"60";
      when x"0299" => bus_data_in <= x"30";
      when x"029a" => bus_data_in <= x"18";
      when x"029b" => bus_data_in <= x"18";
      when x"029c" => bus_data_in <= x"18";
      when x"029d" => bus_data_in <= x"30";
      when x"029e" => bus_data_in <= x"60";
      when x"02a1" => bus_data_in <= x"66";
      when x"02a2" => bus_data_in <= x"3c";
      when x"02a3" => bus_data_in <= x"ff";
      when x"02a4" => bus_data_in <= x"3c";
      when x"02a5" => bus_data_in <= x"66";
      when x"02a9" => bus_data_in <= x"30";
      when x"02aa" => bus_data_in <= x"30";
      when x"02ab" => bus_data_in <= x"fc";
      when x"02ac" => bus_data_in <= x"30";
      when x"02ad" => bus_data_in <= x"30";
      when x"02b5" => bus_data_in <= x"30";
      when x"02b6" => bus_data_in <= x"30";
      when x"02b7" => bus_data_in <= x"60";
      when x"02bb" => bus_data_in <= x"fc";
      when x"02c5" => bus_data_in <= x"30";
      when x"02c6" => bus_data_in <= x"30";
      when x"02c8" => bus_data_in <= x"06";
      when x"02c9" => bus_data_in <= x"0c";
      when x"02ca" => bus_data_in <= x"18";
      when x"02cb" => bus_data_in <= x"30";
      when x"02cc" => bus_data_in <= x"60";
      when x"02cd" => bus_data_in <= x"c0";
      when x"02ce" => bus_data_in <= x"80";
      when x"02d0" => bus_data_in <= x"7c";
      when x"02d1" => bus_data_in <= x"c6";
      when x"02d2" => bus_data_in <= x"ce";
      when x"02d3" => bus_data_in <= x"de";
      when x"02d4" => bus_data_in <= x"f6";
      when x"02d5" => bus_data_in <= x"e6";
      when x"02d6" => bus_data_in <= x"7c";
      when x"02d8" => bus_data_in <= x"30";
      when x"02d9" => bus_data_in <= x"70";
      when x"02da" => bus_data_in <= x"30";
      when x"02db" => bus_data_in <= x"30";
      when x"02dc" => bus_data_in <= x"30";
      when x"02dd" => bus_data_in <= x"30";
      when x"02de" => bus_data_in <= x"fc";
      when x"02e0" => bus_data_in <= x"78";
      when x"02e1" => bus_data_in <= x"cc";
      when x"02e2" => bus_data_in <= x"0c";
      when x"02e3" => bus_data_in <= x"38";
      when x"02e4" => bus_data_in <= x"60";
      when x"02e5" => bus_data_in <= x"cc";
      when x"02e6" => bus_data_in <= x"fc";
      when x"02e8" => bus_data_in <= x"78";
      when x"02e9" => bus_data_in <= x"cc";
      when x"02ea" => bus_data_in <= x"0c";
      when x"02eb" => bus_data_in <= x"38";
      when x"02ec" => bus_data_in <= x"0c";
      when x"02ed" => bus_data_in <= x"cc";
      when x"02ee" => bus_data_in <= x"78";
      when x"02f0" => bus_data_in <= x"1c";
      when x"02f1" => bus_data_in <= x"3c";
      when x"02f2" => bus_data_in <= x"6c";
      when x"02f3" => bus_data_in <= x"cc";
      when x"02f4" => bus_data_in <= x"fe";
      when x"02f5" => bus_data_in <= x"0c";
      when x"02f6" => bus_data_in <= x"1e";
      when x"02f8" => bus_data_in <= x"fc";
      when x"02f9" => bus_data_in <= x"c0";
      when x"02fa" => bus_data_in <= x"f8";
      when x"02fb" => bus_data_in <= x"0c";
      when x"02fc" => bus_data_in <= x"0c";
      when x"02fd" => bus_data_in <= x"cc";
      when x"02fe" => bus_data_in <= x"78";
      when x"0300" => bus_data_in <= x"38";
      when x"0301" => bus_data_in <= x"60";
      when x"0302" => bus_data_in <= x"c0";
      when x"0303" => bus_data_in <= x"f8";
      when x"0304" => bus_data_in <= x"cc";
      when x"0305" => bus_data_in <= x"cc";
      when x"0306" => bus_data_in <= x"78";
      when x"0308" => bus_data_in <= x"fc";
      when x"0309" => bus_data_in <= x"cc";
      when x"030a" => bus_data_in <= x"0c";
      when x"030b" => bus_data_in <= x"18";
      when x"030c" => bus_data_in <= x"30";
      when x"030d" => bus_data_in <= x"30";
      when x"030e" => bus_data_in <= x"30";
      when x"0310" => bus_data_in <= x"78";
      when x"0311" => bus_data_in <= x"cc";
      when x"0312" => bus_data_in <= x"cc";
      when x"0313" => bus_data_in <= x"78";
      when x"0314" => bus_data_in <= x"cc";
      when x"0315" => bus_data_in <= x"cc";
      when x"0316" => bus_data_in <= x"78";
      when x"0318" => bus_data_in <= x"78";
      when x"0319" => bus_data_in <= x"cc";
      when x"031a" => bus_data_in <= x"cc";
      when x"031b" => bus_data_in <= x"7c";
      when x"031c" => bus_data_in <= x"0c";
      when x"031d" => bus_data_in <= x"18";
      when x"031e" => bus_data_in <= x"70";
      when x"0321" => bus_data_in <= x"30";
      when x"0322" => bus_data_in <= x"30";
      when x"0325" => bus_data_in <= x"30";
      when x"0326" => bus_data_in <= x"30";
      when x"0329" => bus_data_in <= x"30";
      when x"032a" => bus_data_in <= x"30";
      when x"032d" => bus_data_in <= x"30";
      when x"032e" => bus_data_in <= x"30";
      when x"032f" => bus_data_in <= x"60";
      when x"0330" => bus_data_in <= x"18";
      when x"0331" => bus_data_in <= x"30";
      when x"0332" => bus_data_in <= x"60";
      when x"0333" => bus_data_in <= x"c0";
      when x"0334" => bus_data_in <= x"60";
      when x"0335" => bus_data_in <= x"30";
      when x"0336" => bus_data_in <= x"18";
      when x"033a" => bus_data_in <= x"fc";
      when x"033d" => bus_data_in <= x"fc";
      when x"0340" => bus_data_in <= x"60";
      when x"0341" => bus_data_in <= x"30";
      when x"0342" => bus_data_in <= x"18";
      when x"0343" => bus_data_in <= x"0c";
      when x"0344" => bus_data_in <= x"18";
      when x"0345" => bus_data_in <= x"30";
      when x"0346" => bus_data_in <= x"60";
      when x"0348" => bus_data_in <= x"78";
      when x"0349" => bus_data_in <= x"cc";
      when x"034a" => bus_data_in <= x"0c";
      when x"034b" => bus_data_in <= x"18";
      when x"034c" => bus_data_in <= x"30";
      when x"034e" => bus_data_in <= x"30";
      when x"0350" => bus_data_in <= x"7c";
      when x"0351" => bus_data_in <= x"c6";
      when x"0352" => bus_data_in <= x"de";
      when x"0353" => bus_data_in <= x"de";
      when x"0354" => bus_data_in <= x"de";
      when x"0355" => bus_data_in <= x"c0";
      when x"0356" => bus_data_in <= x"78";
      when x"0358" => bus_data_in <= x"30";
      when x"0359" => bus_data_in <= x"78";
      when x"035a" => bus_data_in <= x"cc";
      when x"035b" => bus_data_in <= x"cc";
      when x"035c" => bus_data_in <= x"fc";
      when x"035d" => bus_data_in <= x"cc";
      when x"035e" => bus_data_in <= x"cc";
      when x"0360" => bus_data_in <= x"fc";
      when x"0361" => bus_data_in <= x"66";
      when x"0362" => bus_data_in <= x"66";
      when x"0363" => bus_data_in <= x"7c";
      when x"0364" => bus_data_in <= x"66";
      when x"0365" => bus_data_in <= x"66";
      when x"0366" => bus_data_in <= x"fc";
      when x"0368" => bus_data_in <= x"3c";
      when x"0369" => bus_data_in <= x"66";
      when x"036a" => bus_data_in <= x"c0";
      when x"036b" => bus_data_in <= x"c0";
      when x"036c" => bus_data_in <= x"c0";
      when x"036d" => bus_data_in <= x"66";
      when x"036e" => bus_data_in <= x"3c";
      when x"0370" => bus_data_in <= x"f8";
      when x"0371" => bus_data_in <= x"6c";
      when x"0372" => bus_data_in <= x"66";
      when x"0373" => bus_data_in <= x"66";
      when x"0374" => bus_data_in <= x"66";
      when x"0375" => bus_data_in <= x"6c";
      when x"0376" => bus_data_in <= x"f8";
      when x"0378" => bus_data_in <= x"7e";
      when x"0379" => bus_data_in <= x"60";
      when x"037a" => bus_data_in <= x"60";
      when x"037b" => bus_data_in <= x"78";
      when x"037c" => bus_data_in <= x"60";
      when x"037d" => bus_data_in <= x"60";
      when x"037e" => bus_data_in <= x"7e";
      when x"0380" => bus_data_in <= x"7e";
      when x"0381" => bus_data_in <= x"60";
      when x"0382" => bus_data_in <= x"60";
      when x"0383" => bus_data_in <= x"78";
      when x"0384" => bus_data_in <= x"60";
      when x"0385" => bus_data_in <= x"60";
      when x"0386" => bus_data_in <= x"60";
      when x"0388" => bus_data_in <= x"3c";
      when x"0389" => bus_data_in <= x"66";
      when x"038a" => bus_data_in <= x"c0";
      when x"038b" => bus_data_in <= x"c0";
      when x"038c" => bus_data_in <= x"ce";
      when x"038d" => bus_data_in <= x"66";
      when x"038e" => bus_data_in <= x"3e";
      when x"0390" => bus_data_in <= x"cc";
      when x"0391" => bus_data_in <= x"cc";
      when x"0392" => bus_data_in <= x"cc";
      when x"0393" => bus_data_in <= x"fc";
      when x"0394" => bus_data_in <= x"cc";
      when x"0395" => bus_data_in <= x"cc";
      when x"0396" => bus_data_in <= x"cc";
      when x"0398" => bus_data_in <= x"78";
      when x"0399" => bus_data_in <= x"30";
      when x"039a" => bus_data_in <= x"30";
      when x"039b" => bus_data_in <= x"30";
      when x"039c" => bus_data_in <= x"30";
      when x"039d" => bus_data_in <= x"30";
      when x"039e" => bus_data_in <= x"78";
      when x"03a0" => bus_data_in <= x"1e";
      when x"03a1" => bus_data_in <= x"0c";
      when x"03a2" => bus_data_in <= x"0c";
      when x"03a3" => bus_data_in <= x"0c";
      when x"03a4" => bus_data_in <= x"cc";
      when x"03a5" => bus_data_in <= x"cc";
      when x"03a6" => bus_data_in <= x"78";
      when x"03a8" => bus_data_in <= x"e6";
      when x"03a9" => bus_data_in <= x"66";
      when x"03aa" => bus_data_in <= x"6c";
      when x"03ab" => bus_data_in <= x"78";
      when x"03ac" => bus_data_in <= x"6c";
      when x"03ad" => bus_data_in <= x"66";
      when x"03ae" => bus_data_in <= x"e6";
      when x"03b0" => bus_data_in <= x"60";
      when x"03b1" => bus_data_in <= x"60";
      when x"03b2" => bus_data_in <= x"60";
      when x"03b3" => bus_data_in <= x"60";
      when x"03b4" => bus_data_in <= x"60";
      when x"03b5" => bus_data_in <= x"60";
      when x"03b6" => bus_data_in <= x"7e";
      when x"03b8" => bus_data_in <= x"c6";
      when x"03b9" => bus_data_in <= x"ee";
      when x"03ba" => bus_data_in <= x"fe";
      when x"03bb" => bus_data_in <= x"fe";
      when x"03bc" => bus_data_in <= x"d6";
      when x"03bd" => bus_data_in <= x"c6";
      when x"03be" => bus_data_in <= x"c6";
      when x"03c0" => bus_data_in <= x"c6";
      when x"03c1" => bus_data_in <= x"e6";
      when x"03c2" => bus_data_in <= x"f6";
      when x"03c3" => bus_data_in <= x"de";
      when x"03c4" => bus_data_in <= x"ce";
      when x"03c5" => bus_data_in <= x"c6";
      when x"03c6" => bus_data_in <= x"c6";
      when x"03c8" => bus_data_in <= x"38";
      when x"03c9" => bus_data_in <= x"6c";
      when x"03ca" => bus_data_in <= x"c6";
      when x"03cb" => bus_data_in <= x"c6";
      when x"03cc" => bus_data_in <= x"c6";
      when x"03cd" => bus_data_in <= x"6c";
      when x"03ce" => bus_data_in <= x"38";
      when x"03d0" => bus_data_in <= x"fc";
      when x"03d1" => bus_data_in <= x"66";
      when x"03d2" => bus_data_in <= x"66";
      when x"03d3" => bus_data_in <= x"7c";
      when x"03d4" => bus_data_in <= x"60";
      when x"03d5" => bus_data_in <= x"60";
      when x"03d6" => bus_data_in <= x"f0";
      when x"03d8" => bus_data_in <= x"78";
      when x"03d9" => bus_data_in <= x"cc";
      when x"03da" => bus_data_in <= x"cc";
      when x"03db" => bus_data_in <= x"cc";
      when x"03dc" => bus_data_in <= x"dc";
      when x"03dd" => bus_data_in <= x"78";
      when x"03de" => bus_data_in <= x"1c";
      when x"03e0" => bus_data_in <= x"fc";
      when x"03e1" => bus_data_in <= x"66";
      when x"03e2" => bus_data_in <= x"66";
      when x"03e3" => bus_data_in <= x"7c";
      when x"03e4" => bus_data_in <= x"6c";
      when x"03e5" => bus_data_in <= x"66";
      when x"03e6" => bus_data_in <= x"e6";
      when x"03e8" => bus_data_in <= x"78";
      when x"03e9" => bus_data_in <= x"cc";
      when x"03ea" => bus_data_in <= x"e0";
      when x"03eb" => bus_data_in <= x"78";
      when x"03ec" => bus_data_in <= x"1c";
      when x"03ed" => bus_data_in <= x"cc";
      when x"03ee" => bus_data_in <= x"78";
      when x"03f0" => bus_data_in <= x"fc";
      when x"03f1" => bus_data_in <= x"30";
      when x"03f2" => bus_data_in <= x"30";
      when x"03f3" => bus_data_in <= x"30";
      when x"03f4" => bus_data_in <= x"30";
      when x"03f5" => bus_data_in <= x"30";
      when x"03f6" => bus_data_in <= x"30";
      when x"03f8" => bus_data_in <= x"cc";
      when x"03f9" => bus_data_in <= x"cc";
      when x"03fa" => bus_data_in <= x"cc";
      when x"03fb" => bus_data_in <= x"cc";
      when x"03fc" => bus_data_in <= x"cc";
      when x"03fd" => bus_data_in <= x"cc";
      when x"03fe" => bus_data_in <= x"fc";
      when x"0400" => bus_data_in <= x"cc";
      when x"0401" => bus_data_in <= x"cc";
      when x"0402" => bus_data_in <= x"cc";
      when x"0403" => bus_data_in <= x"cc";
      when x"0404" => bus_data_in <= x"cc";
      when x"0405" => bus_data_in <= x"78";
      when x"0406" => bus_data_in <= x"30";
      when x"0408" => bus_data_in <= x"c6";
      when x"0409" => bus_data_in <= x"c6";
      when x"040a" => bus_data_in <= x"c6";
      when x"040b" => bus_data_in <= x"d6";
      when x"040c" => bus_data_in <= x"fe";
      when x"040d" => bus_data_in <= x"ee";
      when x"040e" => bus_data_in <= x"c6";
      when x"0410" => bus_data_in <= x"c6";
      when x"0411" => bus_data_in <= x"c6";
      when x"0412" => bus_data_in <= x"6c";
      when x"0413" => bus_data_in <= x"38";
      when x"0414" => bus_data_in <= x"38";
      when x"0415" => bus_data_in <= x"6c";
      when x"0416" => bus_data_in <= x"c6";
      when x"0418" => bus_data_in <= x"cc";
      when x"0419" => bus_data_in <= x"cc";
      when x"041a" => bus_data_in <= x"cc";
      when x"041b" => bus_data_in <= x"78";
      when x"041c" => bus_data_in <= x"30";
      when x"041d" => bus_data_in <= x"30";
      when x"041e" => bus_data_in <= x"78";
      when x"0420" => bus_data_in <= x"fe";
      when x"0421" => bus_data_in <= x"06";
      when x"0422" => bus_data_in <= x"0c";
      when x"0423" => bus_data_in <= x"18";
      when x"0424" => bus_data_in <= x"30";
      when x"0425" => bus_data_in <= x"60";
      when x"0426" => bus_data_in <= x"fe";
      when x"0428" => bus_data_in <= x"78";
      when x"0429" => bus_data_in <= x"60";
      when x"042a" => bus_data_in <= x"60";
      when x"042b" => bus_data_in <= x"60";
      when x"042c" => bus_data_in <= x"60";
      when x"042d" => bus_data_in <= x"60";
      when x"042e" => bus_data_in <= x"78";
      when x"0430" => bus_data_in <= x"c0";
      when x"0431" => bus_data_in <= x"60";
      when x"0432" => bus_data_in <= x"30";
      when x"0433" => bus_data_in <= x"18";
      when x"0434" => bus_data_in <= x"0c";
      when x"0435" => bus_data_in <= x"06";
      when x"0436" => bus_data_in <= x"02";
      when x"0438" => bus_data_in <= x"78";
      when x"0439" => bus_data_in <= x"18";
      when x"043a" => bus_data_in <= x"18";
      when x"043b" => bus_data_in <= x"18";
      when x"043c" => bus_data_in <= x"18";
      when x"043d" => bus_data_in <= x"18";
      when x"043e" => bus_data_in <= x"78";
      when x"0440" => bus_data_in <= x"10";
      when x"0441" => bus_data_in <= x"38";
      when x"0442" => bus_data_in <= x"6c";
      when x"0443" => bus_data_in <= x"c6";
      when x"044f" => bus_data_in <= x"ff";
      when x"0450" => bus_data_in <= x"30";
      when x"0451" => bus_data_in <= x"30";
      when x"0452" => bus_data_in <= x"18";
      when x"045a" => bus_data_in <= x"78";
      when x"045b" => bus_data_in <= x"0c";
      when x"045c" => bus_data_in <= x"7c";
      when x"045d" => bus_data_in <= x"cc";
      when x"045e" => bus_data_in <= x"76";
      when x"0460" => bus_data_in <= x"e0";
      when x"0461" => bus_data_in <= x"60";
      when x"0462" => bus_data_in <= x"60";
      when x"0463" => bus_data_in <= x"7c";
      when x"0464" => bus_data_in <= x"66";
      when x"0465" => bus_data_in <= x"66";
      when x"0466" => bus_data_in <= x"dc";
      when x"046a" => bus_data_in <= x"78";
      when x"046b" => bus_data_in <= x"cc";
      when x"046c" => bus_data_in <= x"c0";
      when x"046d" => bus_data_in <= x"cc";
      when x"046e" => bus_data_in <= x"78";
      when x"0470" => bus_data_in <= x"1c";
      when x"0471" => bus_data_in <= x"0c";
      when x"0472" => bus_data_in <= x"0c";
      when x"0473" => bus_data_in <= x"7c";
      when x"0474" => bus_data_in <= x"cc";
      when x"0475" => bus_data_in <= x"cc";
      when x"0476" => bus_data_in <= x"76";
      when x"047a" => bus_data_in <= x"78";
      when x"047b" => bus_data_in <= x"cc";
      when x"047c" => bus_data_in <= x"fc";
      when x"047d" => bus_data_in <= x"c0";
      when x"047e" => bus_data_in <= x"78";
      when x"0480" => bus_data_in <= x"38";
      when x"0481" => bus_data_in <= x"6c";
      when x"0482" => bus_data_in <= x"60";
      when x"0483" => bus_data_in <= x"f0";
      when x"0484" => bus_data_in <= x"60";
      when x"0485" => bus_data_in <= x"60";
      when x"0486" => bus_data_in <= x"f0";
      when x"048a" => bus_data_in <= x"76";
      when x"048b" => bus_data_in <= x"cc";
      when x"048c" => bus_data_in <= x"cc";
      when x"048d" => bus_data_in <= x"7c";
      when x"048e" => bus_data_in <= x"0c";
      when x"048f" => bus_data_in <= x"f8";
      when x"0490" => bus_data_in <= x"e0";
      when x"0491" => bus_data_in <= x"60";
      when x"0492" => bus_data_in <= x"6c";
      when x"0493" => bus_data_in <= x"76";
      when x"0494" => bus_data_in <= x"66";
      when x"0495" => bus_data_in <= x"66";
      when x"0496" => bus_data_in <= x"e6";
      when x"0498" => bus_data_in <= x"30";
      when x"049a" => bus_data_in <= x"70";
      when x"049b" => bus_data_in <= x"30";
      when x"049c" => bus_data_in <= x"30";
      when x"049d" => bus_data_in <= x"30";
      when x"049e" => bus_data_in <= x"78";
      when x"04a0" => bus_data_in <= x"0c";
      when x"04a2" => bus_data_in <= x"0c";
      when x"04a3" => bus_data_in <= x"0c";
      when x"04a4" => bus_data_in <= x"0c";
      when x"04a5" => bus_data_in <= x"cc";
      when x"04a6" => bus_data_in <= x"cc";
      when x"04a7" => bus_data_in <= x"78";
      when x"04a8" => bus_data_in <= x"e0";
      when x"04a9" => bus_data_in <= x"60";
      when x"04aa" => bus_data_in <= x"66";
      when x"04ab" => bus_data_in <= x"6c";
      when x"04ac" => bus_data_in <= x"78";
      when x"04ad" => bus_data_in <= x"6c";
      when x"04ae" => bus_data_in <= x"e6";
      when x"04b0" => bus_data_in <= x"70";
      when x"04b1" => bus_data_in <= x"30";
      when x"04b2" => bus_data_in <= x"30";
      when x"04b3" => bus_data_in <= x"30";
      when x"04b4" => bus_data_in <= x"30";
      when x"04b5" => bus_data_in <= x"30";
      when x"04b6" => bus_data_in <= x"78";
      when x"04ba" => bus_data_in <= x"cc";
      when x"04bb" => bus_data_in <= x"fe";
      when x"04bc" => bus_data_in <= x"fe";
      when x"04bd" => bus_data_in <= x"d6";
      when x"04be" => bus_data_in <= x"c6";
      when x"04c2" => bus_data_in <= x"f8";
      when x"04c3" => bus_data_in <= x"cc";
      when x"04c4" => bus_data_in <= x"cc";
      when x"04c5" => bus_data_in <= x"cc";
      when x"04c6" => bus_data_in <= x"cc";
      when x"04ca" => bus_data_in <= x"78";
      when x"04cb" => bus_data_in <= x"cc";
      when x"04cc" => bus_data_in <= x"cc";
      when x"04cd" => bus_data_in <= x"cc";
      when x"04ce" => bus_data_in <= x"78";
      when x"04d2" => bus_data_in <= x"dc";
      when x"04d3" => bus_data_in <= x"66";
      when x"04d4" => bus_data_in <= x"66";
      when x"04d5" => bus_data_in <= x"7c";
      when x"04d6" => bus_data_in <= x"60";
      when x"04d7" => bus_data_in <= x"f0";
      when x"04da" => bus_data_in <= x"76";
      when x"04db" => bus_data_in <= x"cc";
      when x"04dc" => bus_data_in <= x"cc";
      when x"04dd" => bus_data_in <= x"7c";
      when x"04de" => bus_data_in <= x"0c";
      when x"04df" => bus_data_in <= x"1e";
      when x"04e2" => bus_data_in <= x"dc";
      when x"04e3" => bus_data_in <= x"76";
      when x"04e4" => bus_data_in <= x"66";
      when x"04e5" => bus_data_in <= x"60";
      when x"04e6" => bus_data_in <= x"f0";
      when x"04ea" => bus_data_in <= x"7c";
      when x"04eb" => bus_data_in <= x"c0";
      when x"04ec" => bus_data_in <= x"78";
      when x"04ed" => bus_data_in <= x"0c";
      when x"04ee" => bus_data_in <= x"f8";
      when x"04f0" => bus_data_in <= x"10";
      when x"04f1" => bus_data_in <= x"30";
      when x"04f2" => bus_data_in <= x"7c";
      when x"04f3" => bus_data_in <= x"30";
      when x"04f4" => bus_data_in <= x"30";
      when x"04f5" => bus_data_in <= x"34";
      when x"04f6" => bus_data_in <= x"18";
      when x"04fa" => bus_data_in <= x"cc";
      when x"04fb" => bus_data_in <= x"cc";
      when x"04fc" => bus_data_in <= x"cc";
      when x"04fd" => bus_data_in <= x"cc";
      when x"04fe" => bus_data_in <= x"76";
      when x"0502" => bus_data_in <= x"cc";
      when x"0503" => bus_data_in <= x"cc";
      when x"0504" => bus_data_in <= x"cc";
      when x"0505" => bus_data_in <= x"78";
      when x"0506" => bus_data_in <= x"30";
      when x"050a" => bus_data_in <= x"c6";
      when x"050b" => bus_data_in <= x"d6";
      when x"050c" => bus_data_in <= x"fe";
      when x"050d" => bus_data_in <= x"fe";
      when x"050e" => bus_data_in <= x"6c";
      when x"0512" => bus_data_in <= x"c6";
      when x"0513" => bus_data_in <= x"6c";
      when x"0514" => bus_data_in <= x"38";
      when x"0515" => bus_data_in <= x"6c";
      when x"0516" => bus_data_in <= x"c6";
      when x"051a" => bus_data_in <= x"cc";
      when x"051b" => bus_data_in <= x"cc";
      when x"051c" => bus_data_in <= x"cc";
      when x"051d" => bus_data_in <= x"7c";
      when x"051e" => bus_data_in <= x"0c";
      when x"051f" => bus_data_in <= x"f8";
      when x"0522" => bus_data_in <= x"fc";
      when x"0523" => bus_data_in <= x"98";
      when x"0524" => bus_data_in <= x"30";
      when x"0525" => bus_data_in <= x"64";
      when x"0526" => bus_data_in <= x"fc";
      when x"0528" => bus_data_in <= x"1c";
      when x"0529" => bus_data_in <= x"30";
      when x"052a" => bus_data_in <= x"30";
      when x"052b" => bus_data_in <= x"e0";
      when x"052c" => bus_data_in <= x"30";
      when x"052d" => bus_data_in <= x"30";
      when x"052e" => bus_data_in <= x"1c";
      when x"0530" => bus_data_in <= x"18";
      when x"0531" => bus_data_in <= x"18";
      when x"0532" => bus_data_in <= x"18";
      when x"0534" => bus_data_in <= x"18";
      when x"0535" => bus_data_in <= x"18";
      when x"0536" => bus_data_in <= x"18";
      when x"0538" => bus_data_in <= x"e0";
      when x"0539" => bus_data_in <= x"30";
      when x"053a" => bus_data_in <= x"30";
      when x"053b" => bus_data_in <= x"1c";
      when x"053c" => bus_data_in <= x"30";
      when x"053d" => bus_data_in <= x"30";
      when x"053e" => bus_data_in <= x"e0";
      when x"0540" => bus_data_in <= x"76";
      when x"0541" => bus_data_in <= x"dc";
      when x"0549" => bus_data_in <= x"10";
      when x"054a" => bus_data_in <= x"38";
      when x"054b" => bus_data_in <= x"6c";
      when x"054c" => bus_data_in <= x"c6";
      when x"054d" => bus_data_in <= x"fe";
      when x"0550" => bus_data_in <= x"3c";
      when x"0551" => bus_data_in <= x"66";
      when x"0552" => bus_data_in <= x"c0";
      when x"0553" => bus_data_in <= x"c0";
      when x"0554" => bus_data_in <= x"66";
      when x"0555" => bus_data_in <= x"3c";
      when x"0556" => bus_data_in <= x"08";
      when x"0557" => bus_data_in <= x"18";
      when x"0558" => bus_data_in <= x"28";
      when x"055a" => bus_data_in <= x"cc";
      when x"055b" => bus_data_in <= x"cc";
      when x"055c" => bus_data_in <= x"cc";
      when x"055d" => bus_data_in <= x"cc";
      when x"055e" => bus_data_in <= x"76";
      when x"0560" => bus_data_in <= x"08";
      when x"0561" => bus_data_in <= x"10";
      when x"0562" => bus_data_in <= x"78";
      when x"0563" => bus_data_in <= x"cc";
      when x"0564" => bus_data_in <= x"fc";
      when x"0565" => bus_data_in <= x"c0";
      when x"0566" => bus_data_in <= x"78";
      when x"0568" => bus_data_in <= x"10";
      when x"0569" => bus_data_in <= x"28";
      when x"056a" => bus_data_in <= x"78";
      when x"056b" => bus_data_in <= x"0c";
      when x"056c" => bus_data_in <= x"7c";
      when x"056d" => bus_data_in <= x"cc";
      when x"056e" => bus_data_in <= x"76";
      when x"0570" => bus_data_in <= x"28";
      when x"0572" => bus_data_in <= x"78";
      when x"0573" => bus_data_in <= x"0c";
      when x"0574" => bus_data_in <= x"7c";
      when x"0575" => bus_data_in <= x"cc";
      when x"0576" => bus_data_in <= x"76";
      when x"0578" => bus_data_in <= x"20";
      when x"0579" => bus_data_in <= x"10";
      when x"057a" => bus_data_in <= x"78";
      when x"057b" => bus_data_in <= x"0c";
      when x"057c" => bus_data_in <= x"7c";
      when x"057d" => bus_data_in <= x"cc";
      when x"057e" => bus_data_in <= x"76";
      when x"0580" => bus_data_in <= x"18";
      when x"0581" => bus_data_in <= x"18";
      when x"0582" => bus_data_in <= x"78";
      when x"0583" => bus_data_in <= x"0c";
      when x"0584" => bus_data_in <= x"7c";
      when x"0585" => bus_data_in <= x"cc";
      when x"0586" => bus_data_in <= x"76";
      when x"0589" => bus_data_in <= x"78";
      when x"058a" => bus_data_in <= x"cc";
      when x"058b" => bus_data_in <= x"c0";
      when x"058c" => bus_data_in <= x"cc";
      when x"058d" => bus_data_in <= x"78";
      when x"058e" => bus_data_in <= x"10";
      when x"058f" => bus_data_in <= x"30";
      when x"0590" => bus_data_in <= x"10";
      when x"0591" => bus_data_in <= x"28";
      when x"0592" => bus_data_in <= x"78";
      when x"0593" => bus_data_in <= x"cc";
      when x"0594" => bus_data_in <= x"fc";
      when x"0595" => bus_data_in <= x"c0";
      when x"0596" => bus_data_in <= x"78";
      when x"0598" => bus_data_in <= x"28";
      when x"059a" => bus_data_in <= x"78";
      when x"059b" => bus_data_in <= x"cc";
      when x"059c" => bus_data_in <= x"fc";
      when x"059d" => bus_data_in <= x"c0";
      when x"059e" => bus_data_in <= x"78";
      when x"05a0" => bus_data_in <= x"20";
      when x"05a1" => bus_data_in <= x"10";
      when x"05a2" => bus_data_in <= x"78";
      when x"05a3" => bus_data_in <= x"cc";
      when x"05a4" => bus_data_in <= x"fc";
      when x"05a5" => bus_data_in <= x"c0";
      when x"05a6" => bus_data_in <= x"78";
      when x"05a8" => bus_data_in <= x"28";
      when x"05aa" => bus_data_in <= x"70";
      when x"05ab" => bus_data_in <= x"30";
      when x"05ac" => bus_data_in <= x"30";
      when x"05ad" => bus_data_in <= x"30";
      when x"05ae" => bus_data_in <= x"78";
      when x"05b0" => bus_data_in <= x"10";
      when x"05b1" => bus_data_in <= x"28";
      when x"05b2" => bus_data_in <= x"70";
      when x"05b3" => bus_data_in <= x"30";
      when x"05b4" => bus_data_in <= x"30";
      when x"05b5" => bus_data_in <= x"30";
      when x"05b6" => bus_data_in <= x"78";
      when x"05b8" => bus_data_in <= x"10";
      when x"05b9" => bus_data_in <= x"08";
      when x"05ba" => bus_data_in <= x"70";
      when x"05bb" => bus_data_in <= x"30";
      when x"05bc" => bus_data_in <= x"30";
      when x"05bd" => bus_data_in <= x"30";
      when x"05be" => bus_data_in <= x"78";
      when x"05c0" => bus_data_in <= x"28";
      when x"05c1" => bus_data_in <= x"30";
      when x"05c2" => bus_data_in <= x"78";
      when x"05c3" => bus_data_in <= x"cc";
      when x"05c4" => bus_data_in <= x"fc";
      when x"05c5" => bus_data_in <= x"cc";
      when x"05c6" => bus_data_in <= x"cc";
      when x"05c8" => bus_data_in <= x"30";
      when x"05c9" => bus_data_in <= x"48";
      when x"05ca" => bus_data_in <= x"30";
      when x"05cb" => bus_data_in <= x"cc";
      when x"05cc" => bus_data_in <= x"fc";
      when x"05cd" => bus_data_in <= x"cc";
      when x"05ce" => bus_data_in <= x"cc";
      when x"05d0" => bus_data_in <= x"08";
      when x"05d1" => bus_data_in <= x"10";
      when x"05d2" => bus_data_in <= x"7e";
      when x"05d3" => bus_data_in <= x"60";
      when x"05d4" => bus_data_in <= x"78";
      when x"05d5" => bus_data_in <= x"60";
      when x"05d6" => bus_data_in <= x"7e";
      when x"05da" => bus_data_in <= x"6c";
      when x"05db" => bus_data_in <= x"12";
      when x"05dc" => bus_data_in <= x"7e";
      when x"05dd" => bus_data_in <= x"90";
      when x"05de" => bus_data_in <= x"7e";
      when x"05e0" => bus_data_in <= x"3e";
      when x"05e1" => bus_data_in <= x"50";
      when x"05e2" => bus_data_in <= x"90";
      when x"05e3" => bus_data_in <= x"9c";
      when x"05e4" => bus_data_in <= x"f0";
      when x"05e5" => bus_data_in <= x"90";
      when x"05e6" => bus_data_in <= x"9e";
      when x"05e8" => bus_data_in <= x"10";
      when x"05e9" => bus_data_in <= x"28";
      when x"05ea" => bus_data_in <= x"78";
      when x"05eb" => bus_data_in <= x"cc";
      when x"05ec" => bus_data_in <= x"cc";
      when x"05ed" => bus_data_in <= x"cc";
      when x"05ee" => bus_data_in <= x"78";
      when x"05f0" => bus_data_in <= x"28";
      when x"05f2" => bus_data_in <= x"78";
      when x"05f3" => bus_data_in <= x"cc";
      when x"05f4" => bus_data_in <= x"cc";
      when x"05f5" => bus_data_in <= x"cc";
      when x"05f6" => bus_data_in <= x"78";
      when x"05f8" => bus_data_in <= x"20";
      when x"05f9" => bus_data_in <= x"10";
      when x"05fa" => bus_data_in <= x"78";
      when x"05fb" => bus_data_in <= x"cc";
      when x"05fc" => bus_data_in <= x"cc";
      when x"05fd" => bus_data_in <= x"cc";
      when x"05fe" => bus_data_in <= x"78";
      when x"0600" => bus_data_in <= x"10";
      when x"0601" => bus_data_in <= x"28";
      when x"0602" => bus_data_in <= x"cc";
      when x"0603" => bus_data_in <= x"cc";
      when x"0604" => bus_data_in <= x"cc";
      when x"0605" => bus_data_in <= x"cc";
      when x"0606" => bus_data_in <= x"76";
      when x"0608" => bus_data_in <= x"20";
      when x"0609" => bus_data_in <= x"10";
      when x"060a" => bus_data_in <= x"cc";
      when x"060b" => bus_data_in <= x"cc";
      when x"060c" => bus_data_in <= x"cc";
      when x"060d" => bus_data_in <= x"cc";
      when x"060e" => bus_data_in <= x"76";
      when x"0610" => bus_data_in <= x"28";
      when x"0612" => bus_data_in <= x"cc";
      when x"0613" => bus_data_in <= x"cc";
      when x"0614" => bus_data_in <= x"cc";
      when x"0615" => bus_data_in <= x"7c";
      when x"0616" => bus_data_in <= x"0c";
      when x"0617" => bus_data_in <= x"f8";
      when x"0618" => bus_data_in <= x"28";
      when x"0619" => bus_data_in <= x"7c";
      when x"061a" => bus_data_in <= x"c6";
      when x"061b" => bus_data_in <= x"c6";
      when x"061c" => bus_data_in <= x"c6";
      when x"061d" => bus_data_in <= x"c6";
      when x"061e" => bus_data_in <= x"7c";
      when x"0620" => bus_data_in <= x"28";
      when x"0621" => bus_data_in <= x"c6";
      when x"0622" => bus_data_in <= x"c6";
      when x"0623" => bus_data_in <= x"c6";
      when x"0624" => bus_data_in <= x"c6";
      when x"0625" => bus_data_in <= x"c6";
      when x"0626" => bus_data_in <= x"7c";
      when x"0629" => bus_data_in <= x"10";
      when x"062a" => bus_data_in <= x"78";
      when x"062b" => bus_data_in <= x"cc";
      when x"062c" => bus_data_in <= x"c0";
      when x"062d" => bus_data_in <= x"cc";
      when x"062e" => bus_data_in <= x"78";
      when x"062f" => bus_data_in <= x"10";
      when x"0630" => bus_data_in <= x"38";
      when x"0631" => bus_data_in <= x"44";
      when x"0632" => bus_data_in <= x"40";
      when x"0633" => bus_data_in <= x"f0";
      when x"0634" => bus_data_in <= x"40";
      when x"0635" => bus_data_in <= x"40";
      when x"0636" => bus_data_in <= x"fe";
      when x"0638" => bus_data_in <= x"c3";
      when x"0639" => bus_data_in <= x"66";
      when x"063a" => bus_data_in <= x"3c";
      when x"063b" => bus_data_in <= x"7e";
      when x"063c" => bus_data_in <= x"18";
      when x"063d" => bus_data_in <= x"7e";
      when x"063e" => bus_data_in <= x"18";
      when x"0640" => bus_data_in <= x"fc";
      when x"0641" => bus_data_in <= x"66";
      when x"0642" => bus_data_in <= x"66";
      when x"0643" => bus_data_in <= x"7c";
      when x"0644" => bus_data_in <= x"60";
      when x"0645" => bus_data_in <= x"60";
      when x"0646" => bus_data_in <= x"f0";
      when x"0648" => bus_data_in <= x"1c";
      when x"0649" => bus_data_in <= x"30";
      when x"064a" => bus_data_in <= x"fc";
      when x"064b" => bus_data_in <= x"30";
      when x"064c" => bus_data_in <= x"30";
      when x"064d" => bus_data_in <= x"30";
      when x"064e" => bus_data_in <= x"30";
      when x"064f" => bus_data_in <= x"e0";
      when x"0650" => bus_data_in <= x"08";
      when x"0651" => bus_data_in <= x"10";
      when x"0652" => bus_data_in <= x"78";
      when x"0653" => bus_data_in <= x"0c";
      when x"0654" => bus_data_in <= x"7c";
      when x"0655" => bus_data_in <= x"cc";
      when x"0656" => bus_data_in <= x"76";
      when x"0658" => bus_data_in <= x"10";
      when x"0659" => bus_data_in <= x"20";
      when x"065a" => bus_data_in <= x"70";
      when x"065b" => bus_data_in <= x"30";
      when x"065c" => bus_data_in <= x"30";
      when x"065d" => bus_data_in <= x"30";
      when x"065e" => bus_data_in <= x"78";
      when x"0660" => bus_data_in <= x"10";
      when x"0661" => bus_data_in <= x"20";
      when x"0662" => bus_data_in <= x"78";
      when x"0663" => bus_data_in <= x"cc";
      when x"0664" => bus_data_in <= x"cc";
      when x"0665" => bus_data_in <= x"cc";
      when x"0666" => bus_data_in <= x"78";
      when x"0668" => bus_data_in <= x"10";
      when x"0669" => bus_data_in <= x"20";
      when x"066a" => bus_data_in <= x"cc";
      when x"066b" => bus_data_in <= x"cc";
      when x"066c" => bus_data_in <= x"cc";
      when x"066d" => bus_data_in <= x"cc";
      when x"066e" => bus_data_in <= x"76";
      when x"0670" => bus_data_in <= x"32";
      when x"0671" => bus_data_in <= x"4c";
      when x"0672" => bus_data_in <= x"f8";
      when x"0673" => bus_data_in <= x"cc";
      when x"0674" => bus_data_in <= x"cc";
      when x"0675" => bus_data_in <= x"cc";
      when x"0676" => bus_data_in <= x"cc";
      when x"0678" => bus_data_in <= x"32";
      when x"0679" => bus_data_in <= x"4c";
      when x"067a" => bus_data_in <= x"c6";
      when x"067b" => bus_data_in <= x"e6";
      when x"067c" => bus_data_in <= x"d6";
      when x"067d" => bus_data_in <= x"ce";
      when x"067e" => bus_data_in <= x"c6";
      when x"0681" => bus_data_in <= x"38";
      when x"0682" => bus_data_in <= x"0c";
      when x"0683" => bus_data_in <= x"3c";
      when x"0684" => bus_data_in <= x"6c";
      when x"0685" => bus_data_in <= x"36";
      when x"0689" => bus_data_in <= x"38";
      when x"068a" => bus_data_in <= x"44";
      when x"068b" => bus_data_in <= x"44";
      when x"068c" => bus_data_in <= x"38";
      when x"0690" => bus_data_in <= x"18";
      when x"0692" => bus_data_in <= x"18";
      when x"0693" => bus_data_in <= x"30";
      when x"0694" => bus_data_in <= x"60";
      when x"0695" => bus_data_in <= x"66";
      when x"0696" => bus_data_in <= x"3c";
      when x"069a" => bus_data_in <= x"fe";
      when x"069b" => bus_data_in <= x"80";
      when x"069c" => bus_data_in <= x"80";
      when x"06a2" => bus_data_in <= x"fe";
      when x"06a3" => bus_data_in <= x"02";
      when x"06a4" => bus_data_in <= x"02";
      when x"06a8" => bus_data_in <= x"42";
      when x"06a9" => bus_data_in <= x"44";
      when x"06aa" => bus_data_in <= x"48";
      when x"06ab" => bus_data_in <= x"56";
      when x"06ac" => bus_data_in <= x"29";
      when x"06ad" => bus_data_in <= x"46";
      when x"06ae" => bus_data_in <= x"88";
      when x"06af" => bus_data_in <= x"1f";
      when x"06b0" => bus_data_in <= x"42";
      when x"06b1" => bus_data_in <= x"44";
      when x"06b2" => bus_data_in <= x"48";
      when x"06b3" => bus_data_in <= x"56";
      when x"06b4" => bus_data_in <= x"2a";
      when x"06b5" => bus_data_in <= x"5f";
      when x"06b6" => bus_data_in <= x"82";
      when x"06b7" => bus_data_in <= x"07";
      when x"06b8" => bus_data_in <= x"30";
      when x"06ba" => bus_data_in <= x"30";
      when x"06bb" => bus_data_in <= x"30";
      when x"06bc" => bus_data_in <= x"30";
      when x"06bd" => bus_data_in <= x"30";
      when x"06be" => bus_data_in <= x"30";
      when x"06c1" => bus_data_in <= x"24";
      when x"06c2" => bus_data_in <= x"48";
      when x"06c3" => bus_data_in <= x"90";
      when x"06c4" => bus_data_in <= x"48";
      when x"06c5" => bus_data_in <= x"24";
      when x"06c9" => bus_data_in <= x"48";
      when x"06ca" => bus_data_in <= x"24";
      when x"06cb" => bus_data_in <= x"12";
      when x"06cc" => bus_data_in <= x"24";
      when x"06cd" => bus_data_in <= x"48";
      when x"06d0" => bus_data_in <= x"88";
      when x"06d1" => bus_data_in <= x"22";
      when x"06d2" => bus_data_in <= x"88";
      when x"06d3" => bus_data_in <= x"22";
      when x"06d4" => bus_data_in <= x"88";
      when x"06d6" => bus_data_in <= x"88";
      when x"06d7" => bus_data_in <= x"22";
      when x"06d8" => bus_data_in <= x"aa";
      when x"06d9" => bus_data_in <= x"55";
      when x"06da" => bus_data_in <= x"aa";
      when x"06db" => bus_data_in <= x"55";
      when x"06dc" => bus_data_in <= x"aa";
      when x"06de" => bus_data_in <= x"aa";
      when x"06df" => bus_data_in <= x"55";
      when x"06e0" => bus_data_in <= x"77";
      when x"06e1" => bus_data_in <= x"dd";
      when x"06e2" => bus_data_in <= x"77";
      when x"06e3" => bus_data_in <= x"dd";
      when x"06e4" => bus_data_in <= x"77";
      when x"06e5" => bus_data_in <= x"ff";
      when x"06e6" => bus_data_in <= x"77";
      when x"06e7" => bus_data_in <= x"dd";
      when x"06e8" => bus_data_in <= x"10";
      when x"06e9" => bus_data_in <= x"10";
      when x"06ea" => bus_data_in <= x"10";
      when x"06eb" => bus_data_in <= x"10";
      when x"06ec" => bus_data_in <= x"10";
      when x"06ed" => bus_data_in <= x"10";
      when x"06ee" => bus_data_in <= x"10";
      when x"06ef" => bus_data_in <= x"10";
      when x"06f0" => bus_data_in <= x"10";
      when x"06f1" => bus_data_in <= x"10";
      when x"06f2" => bus_data_in <= x"10";
      when x"06f3" => bus_data_in <= x"f0";
      when x"06f4" => bus_data_in <= x"10";
      when x"06f5" => bus_data_in <= x"10";
      when x"06f6" => bus_data_in <= x"10";
      when x"06f7" => bus_data_in <= x"10";
      when x"06f8" => bus_data_in <= x"10";
      when x"06f9" => bus_data_in <= x"10";
      when x"06fa" => bus_data_in <= x"f0";
      when x"06fb" => bus_data_in <= x"10";
      when x"06fc" => bus_data_in <= x"f0";
      when x"06fd" => bus_data_in <= x"10";
      when x"06fe" => bus_data_in <= x"10";
      when x"06ff" => bus_data_in <= x"10";
      when x"0700" => bus_data_in <= x"28";
      when x"0701" => bus_data_in <= x"28";
      when x"0702" => bus_data_in <= x"28";
      when x"0703" => bus_data_in <= x"e8";
      when x"0704" => bus_data_in <= x"28";
      when x"0705" => bus_data_in <= x"28";
      when x"0706" => bus_data_in <= x"28";
      when x"0707" => bus_data_in <= x"28";
      when x"070b" => bus_data_in <= x"f8";
      when x"070c" => bus_data_in <= x"28";
      when x"070d" => bus_data_in <= x"28";
      when x"070e" => bus_data_in <= x"28";
      when x"070f" => bus_data_in <= x"28";
      when x"0712" => bus_data_in <= x"f0";
      when x"0713" => bus_data_in <= x"10";
      when x"0714" => bus_data_in <= x"f0";
      when x"0715" => bus_data_in <= x"10";
      when x"0716" => bus_data_in <= x"10";
      when x"0717" => bus_data_in <= x"10";
      when x"0718" => bus_data_in <= x"28";
      when x"0719" => bus_data_in <= x"28";
      when x"071a" => bus_data_in <= x"e8";
      when x"071b" => bus_data_in <= x"08";
      when x"071c" => bus_data_in <= x"e8";
      when x"071d" => bus_data_in <= x"28";
      when x"071e" => bus_data_in <= x"28";
      when x"071f" => bus_data_in <= x"28";
      when x"0720" => bus_data_in <= x"28";
      when x"0721" => bus_data_in <= x"28";
      when x"0722" => bus_data_in <= x"28";
      when x"0723" => bus_data_in <= x"28";
      when x"0724" => bus_data_in <= x"28";
      when x"0725" => bus_data_in <= x"28";
      when x"0726" => bus_data_in <= x"28";
      when x"0727" => bus_data_in <= x"28";
      when x"072a" => bus_data_in <= x"f8";
      when x"072b" => bus_data_in <= x"08";
      when x"072c" => bus_data_in <= x"e8";
      when x"072d" => bus_data_in <= x"28";
      when x"072e" => bus_data_in <= x"28";
      when x"072f" => bus_data_in <= x"28";
      when x"0730" => bus_data_in <= x"28";
      when x"0731" => bus_data_in <= x"28";
      when x"0732" => bus_data_in <= x"e8";
      when x"0733" => bus_data_in <= x"08";
      when x"0734" => bus_data_in <= x"f8";
      when x"0738" => bus_data_in <= x"28";
      when x"0739" => bus_data_in <= x"28";
      when x"073a" => bus_data_in <= x"28";
      when x"073b" => bus_data_in <= x"f8";
      when x"0740" => bus_data_in <= x"10";
      when x"0741" => bus_data_in <= x"10";
      when x"0742" => bus_data_in <= x"f0";
      when x"0743" => bus_data_in <= x"10";
      when x"0744" => bus_data_in <= x"f0";
      when x"074b" => bus_data_in <= x"f0";
      when x"074c" => bus_data_in <= x"10";
      when x"074d" => bus_data_in <= x"10";
      when x"074e" => bus_data_in <= x"10";
      when x"074f" => bus_data_in <= x"10";
      when x"0750" => bus_data_in <= x"10";
      when x"0751" => bus_data_in <= x"10";
      when x"0752" => bus_data_in <= x"10";
      when x"0753" => bus_data_in <= x"1f";
      when x"0758" => bus_data_in <= x"10";
      when x"0759" => bus_data_in <= x"10";
      when x"075a" => bus_data_in <= x"10";
      when x"075b" => bus_data_in <= x"ff";
      when x"0763" => bus_data_in <= x"ff";
      when x"0764" => bus_data_in <= x"10";
      when x"0765" => bus_data_in <= x"10";
      when x"0766" => bus_data_in <= x"10";
      when x"0767" => bus_data_in <= x"10";
      when x"0768" => bus_data_in <= x"10";
      when x"0769" => bus_data_in <= x"10";
      when x"076a" => bus_data_in <= x"10";
      when x"076b" => bus_data_in <= x"1f";
      when x"076c" => bus_data_in <= x"10";
      when x"076d" => bus_data_in <= x"10";
      when x"076e" => bus_data_in <= x"10";
      when x"076f" => bus_data_in <= x"10";
      when x"0773" => bus_data_in <= x"ff";
      when x"0778" => bus_data_in <= x"10";
      when x"0779" => bus_data_in <= x"10";
      when x"077a" => bus_data_in <= x"10";
      when x"077b" => bus_data_in <= x"ff";
      when x"077c" => bus_data_in <= x"10";
      when x"077d" => bus_data_in <= x"10";
      when x"077e" => bus_data_in <= x"10";
      when x"077f" => bus_data_in <= x"10";
      when x"0780" => bus_data_in <= x"10";
      when x"0781" => bus_data_in <= x"10";
      when x"0782" => bus_data_in <= x"1f";
      when x"0783" => bus_data_in <= x"10";
      when x"0784" => bus_data_in <= x"1f";
      when x"0785" => bus_data_in <= x"10";
      when x"0786" => bus_data_in <= x"10";
      when x"0787" => bus_data_in <= x"10";
      when x"0788" => bus_data_in <= x"28";
      when x"0789" => bus_data_in <= x"28";
      when x"078a" => bus_data_in <= x"28";
      when x"078b" => bus_data_in <= x"2f";
      when x"078c" => bus_data_in <= x"28";
      when x"078d" => bus_data_in <= x"28";
      when x"078e" => bus_data_in <= x"28";
      when x"078f" => bus_data_in <= x"28";
      when x"0790" => bus_data_in <= x"28";
      when x"0791" => bus_data_in <= x"28";
      when x"0792" => bus_data_in <= x"2f";
      when x"0793" => bus_data_in <= x"20";
      when x"0794" => bus_data_in <= x"3f";
      when x"079a" => bus_data_in <= x"3f";
      when x"079b" => bus_data_in <= x"20";
      when x"079c" => bus_data_in <= x"2f";
      when x"079d" => bus_data_in <= x"28";
      when x"079e" => bus_data_in <= x"28";
      when x"079f" => bus_data_in <= x"28";
      when x"07a0" => bus_data_in <= x"28";
      when x"07a1" => bus_data_in <= x"28";
      when x"07a2" => bus_data_in <= x"ef";
      when x"07a4" => bus_data_in <= x"ff";
      when x"07aa" => bus_data_in <= x"ff";
      when x"07ac" => bus_data_in <= x"ef";
      when x"07ad" => bus_data_in <= x"28";
      when x"07ae" => bus_data_in <= x"28";
      when x"07af" => bus_data_in <= x"28";
      when x"07b0" => bus_data_in <= x"28";
      when x"07b1" => bus_data_in <= x"28";
      when x"07b2" => bus_data_in <= x"2f";
      when x"07b3" => bus_data_in <= x"20";
      when x"07b4" => bus_data_in <= x"2f";
      when x"07b5" => bus_data_in <= x"28";
      when x"07b6" => bus_data_in <= x"28";
      when x"07b7" => bus_data_in <= x"28";
      when x"07ba" => bus_data_in <= x"ff";
      when x"07bc" => bus_data_in <= x"ff";
      when x"07c0" => bus_data_in <= x"28";
      when x"07c1" => bus_data_in <= x"28";
      when x"07c2" => bus_data_in <= x"ef";
      when x"07c4" => bus_data_in <= x"ef";
      when x"07c5" => bus_data_in <= x"28";
      when x"07c6" => bus_data_in <= x"28";
      when x"07c7" => bus_data_in <= x"28";
      when x"07c8" => bus_data_in <= x"10";
      when x"07c9" => bus_data_in <= x"10";
      when x"07ca" => bus_data_in <= x"ff";
      when x"07cc" => bus_data_in <= x"ff";
      when x"07d0" => bus_data_in <= x"28";
      when x"07d1" => bus_data_in <= x"28";
      when x"07d2" => bus_data_in <= x"28";
      when x"07d3" => bus_data_in <= x"ff";
      when x"07da" => bus_data_in <= x"ff";
      when x"07dc" => bus_data_in <= x"ff";
      when x"07dd" => bus_data_in <= x"10";
      when x"07de" => bus_data_in <= x"10";
      when x"07df" => bus_data_in <= x"10";
      when x"07e3" => bus_data_in <= x"ff";
      when x"07e4" => bus_data_in <= x"28";
      when x"07e5" => bus_data_in <= x"28";
      when x"07e6" => bus_data_in <= x"28";
      when x"07e7" => bus_data_in <= x"28";
      when x"07e8" => bus_data_in <= x"28";
      when x"07e9" => bus_data_in <= x"28";
      when x"07ea" => bus_data_in <= x"28";
      when x"07eb" => bus_data_in <= x"3f";
      when x"07f0" => bus_data_in <= x"10";
      when x"07f1" => bus_data_in <= x"10";
      when x"07f2" => bus_data_in <= x"1f";
      when x"07f3" => bus_data_in <= x"10";
      when x"07f4" => bus_data_in <= x"1f";
      when x"07fa" => bus_data_in <= x"1f";
      when x"07fb" => bus_data_in <= x"10";
      when x"07fc" => bus_data_in <= x"1f";
      when x"07fd" => bus_data_in <= x"10";
      when x"07fe" => bus_data_in <= x"10";
      when x"07ff" => bus_data_in <= x"10";
      when x"0803" => bus_data_in <= x"3f";
      when x"0804" => bus_data_in <= x"28";
      when x"0805" => bus_data_in <= x"28";
      when x"0806" => bus_data_in <= x"28";
      when x"0807" => bus_data_in <= x"28";
      when x"0808" => bus_data_in <= x"28";
      when x"0809" => bus_data_in <= x"28";
      when x"080a" => bus_data_in <= x"28";
      when x"080b" => bus_data_in <= x"ff";
      when x"080c" => bus_data_in <= x"28";
      when x"080d" => bus_data_in <= x"28";
      when x"080e" => bus_data_in <= x"28";
      when x"080f" => bus_data_in <= x"28";
      when x"0810" => bus_data_in <= x"10";
      when x"0811" => bus_data_in <= x"10";
      when x"0812" => bus_data_in <= x"ff";
      when x"0813" => bus_data_in <= x"10";
      when x"0814" => bus_data_in <= x"ff";
      when x"0815" => bus_data_in <= x"10";
      when x"0816" => bus_data_in <= x"10";
      when x"0817" => bus_data_in <= x"10";
      when x"0818" => bus_data_in <= x"10";
      when x"0819" => bus_data_in <= x"10";
      when x"081a" => bus_data_in <= x"10";
      when x"081b" => bus_data_in <= x"f0";
      when x"0823" => bus_data_in <= x"1f";
      when x"0824" => bus_data_in <= x"10";
      when x"0825" => bus_data_in <= x"10";
      when x"0826" => bus_data_in <= x"10";
      when x"0827" => bus_data_in <= x"10";
      when x"0828" => bus_data_in <= x"ff";
      when x"0829" => bus_data_in <= x"ff";
      when x"082a" => bus_data_in <= x"ff";
      when x"082b" => bus_data_in <= x"ff";
      when x"082c" => bus_data_in <= x"ff";
      when x"082d" => bus_data_in <= x"ff";
      when x"082e" => bus_data_in <= x"ff";
      when x"082f" => bus_data_in <= x"ff";
      when x"0834" => bus_data_in <= x"ff";
      when x"0835" => bus_data_in <= x"ff";
      when x"0836" => bus_data_in <= x"ff";
      when x"0837" => bus_data_in <= x"ff";
      when x"0838" => bus_data_in <= x"f0";
      when x"0839" => bus_data_in <= x"f0";
      when x"083a" => bus_data_in <= x"f0";
      when x"083b" => bus_data_in <= x"f0";
      when x"083c" => bus_data_in <= x"f0";
      when x"083d" => bus_data_in <= x"f0";
      when x"083e" => bus_data_in <= x"f0";
      when x"083f" => bus_data_in <= x"f0";
      when x"0840" => bus_data_in <= x"0f";
      when x"0841" => bus_data_in <= x"0f";
      when x"0842" => bus_data_in <= x"0f";
      when x"0843" => bus_data_in <= x"0f";
      when x"0844" => bus_data_in <= x"0f";
      when x"0845" => bus_data_in <= x"0f";
      when x"0846" => bus_data_in <= x"0f";
      when x"0847" => bus_data_in <= x"0f";
      when x"0848" => bus_data_in <= x"ff";
      when x"0849" => bus_data_in <= x"ff";
      when x"084a" => bus_data_in <= x"ff";
      when x"084b" => bus_data_in <= x"ff";
      when x"0853" => bus_data_in <= x"72";
      when x"0854" => bus_data_in <= x"8c";
      when x"0855" => bus_data_in <= x"88";
      when x"0856" => bus_data_in <= x"3a";
      when x"0858" => bus_data_in <= x"30";
      when x"0859" => bus_data_in <= x"48";
      when x"085a" => bus_data_in <= x"48";
      when x"085b" => bus_data_in <= x"7c";
      when x"085c" => bus_data_in <= x"42";
      when x"085d" => bus_data_in <= x"42";
      when x"085e" => bus_data_in <= x"dc";
      when x"0862" => bus_data_in <= x"fe";
      when x"0863" => bus_data_in <= x"42";
      when x"0864" => bus_data_in <= x"40";
      when x"0865" => bus_data_in <= x"40";
      when x"0866" => bus_data_in <= x"e0";
      when x"086a" => bus_data_in <= x"fe";
      when x"086b" => bus_data_in <= x"44";
      when x"086c" => bus_data_in <= x"44";
      when x"086d" => bus_data_in <= x"44";
      when x"086e" => bus_data_in <= x"ee";
      when x"0870" => bus_data_in <= x"fe";
      when x"0871" => bus_data_in <= x"42";
      when x"0872" => bus_data_in <= x"20";
      when x"0873" => bus_data_in <= x"10";
      when x"0874" => bus_data_in <= x"20";
      when x"0875" => bus_data_in <= x"42";
      when x"0876" => bus_data_in <= x"fe";
      when x"087b" => bus_data_in <= x"3e";
      when x"087c" => bus_data_in <= x"44";
      when x"087d" => bus_data_in <= x"44";
      when x"087e" => bus_data_in <= x"38";
      when x"0882" => bus_data_in <= x"cc";
      when x"0883" => bus_data_in <= x"44";
      when x"0884" => bus_data_in <= x"44";
      when x"0885" => bus_data_in <= x"44";
      when x"0886" => bus_data_in <= x"7a";
      when x"0887" => bus_data_in <= x"40";
      when x"088a" => bus_data_in <= x"7c";
      when x"088b" => bus_data_in <= x"10";
      when x"088c" => bus_data_in <= x"10";
      when x"088d" => bus_data_in <= x"10";
      when x"088e" => bus_data_in <= x"1c";
      when x"0891" => bus_data_in <= x"10";
      when x"0892" => bus_data_in <= x"7c";
      when x"0893" => bus_data_in <= x"92";
      when x"0894" => bus_data_in <= x"92";
      when x"0895" => bus_data_in <= x"7c";
      when x"0896" => bus_data_in <= x"10";
      when x"089a" => bus_data_in <= x"7c";
      when x"089b" => bus_data_in <= x"82";
      when x"089c" => bus_data_in <= x"ba";
      when x"089d" => bus_data_in <= x"82";
      when x"089e" => bus_data_in <= x"7c";
      when x"08a3" => bus_data_in <= x"7c";
      when x"08a4" => bus_data_in <= x"82";
      when x"08a5" => bus_data_in <= x"82";
      when x"08a6" => bus_data_in <= x"6c";
      when x"08a7" => bus_data_in <= x"28";
      when x"08a8" => bus_data_in <= x"ee";
      when x"08ab" => bus_data_in <= x"7c";
      when x"08ac" => bus_data_in <= x"20";
      when x"08ad" => bus_data_in <= x"38";
      when x"08ae" => bus_data_in <= x"44";
      when x"08af" => bus_data_in <= x"44";
      when x"08b0" => bus_data_in <= x"38";
      when x"08b4" => bus_data_in <= x"6c";
      when x"08b5" => bus_data_in <= x"92";
      when x"08b6" => bus_data_in <= x"92";
      when x"08b7" => bus_data_in <= x"6c";
      when x"08bc" => bus_data_in <= x"4c";
      when x"08bd" => bus_data_in <= x"92";
      when x"08be" => bus_data_in <= x"92";
      when x"08bf" => bus_data_in <= x"7c";
      when x"08c0" => bus_data_in <= x"10";
      when x"08c4" => bus_data_in <= x"3c";
      when x"08c5" => bus_data_in <= x"40";
      when x"08c6" => bus_data_in <= x"30";
      when x"08c7" => bus_data_in <= x"40";
      when x"08c8" => bus_data_in <= x"3c";
      when x"08cc" => bus_data_in <= x"3c";
      when x"08cd" => bus_data_in <= x"42";
      when x"08ce" => bus_data_in <= x"42";
      when x"08cf" => bus_data_in <= x"42";
      when x"08d0" => bus_data_in <= x"42";
      when x"08d3" => bus_data_in <= x"fe";
      when x"08d5" => bus_data_in <= x"fe";
      when x"08d7" => bus_data_in <= x"fe";
      when x"08da" => bus_data_in <= x"10";
      when x"08db" => bus_data_in <= x"10";
      when x"08dc" => bus_data_in <= x"fe";
      when x"08dd" => bus_data_in <= x"10";
      when x"08de" => bus_data_in <= x"10";
      when x"08df" => bus_data_in <= x"fe";
      when x"08e2" => bus_data_in <= x"40";
      when x"08e3" => bus_data_in <= x"10";
      when x"08e4" => bus_data_in <= x"04";
      when x"08e5" => bus_data_in <= x"10";
      when x"08e6" => bus_data_in <= x"40";
      when x"08e7" => bus_data_in <= x"fe";
      when x"08ea" => bus_data_in <= x"04";
      when x"08eb" => bus_data_in <= x"10";
      when x"08ec" => bus_data_in <= x"40";
      when x"08ed" => bus_data_in <= x"10";
      when x"08ee" => bus_data_in <= x"04";
      when x"08ef" => bus_data_in <= x"fe";
      when x"08f2" => bus_data_in <= x"0c";
      when x"08f3" => bus_data_in <= x"10";
      when x"08f4" => bus_data_in <= x"10";
      when x"08f5" => bus_data_in <= x"10";
      when x"08f6" => bus_data_in <= x"10";
      when x"08f7" => bus_data_in <= x"10";
      when x"08f8" => bus_data_in <= x"10";
      when x"08f9" => bus_data_in <= x"10";
      when x"08fa" => bus_data_in <= x"10";
      when x"08fb" => bus_data_in <= x"10";
      when x"08fc" => bus_data_in <= x"10";
      when x"08fd" => bus_data_in <= x"10";
      when x"08fe" => bus_data_in <= x"10";
      when x"08ff" => bus_data_in <= x"10";
      when x"0900" => bus_data_in <= x"10";
      when x"0901" => bus_data_in <= x"60";
      when x"0904" => bus_data_in <= x"10";
      when x"0906" => bus_data_in <= x"fe";
      when x"0908" => bus_data_in <= x"10";
      when x"090b" => bus_data_in <= x"62";
      when x"090c" => bus_data_in <= x"9c";
      when x"090e" => bus_data_in <= x"62";
      when x"090f" => bus_data_in <= x"9c";
      when x"0912" => bus_data_in <= x"30";
      when x"0913" => bus_data_in <= x"48";
      when x"0914" => bus_data_in <= x"48";
      when x"0915" => bus_data_in <= x"30";
      when x"091d" => bus_data_in <= x"30";
      when x"091e" => bus_data_in <= x"30";
      when x"0926" => bus_data_in <= x"08";
      when x"092a" => bus_data_in <= x"01";
      when x"092b" => bus_data_in <= x"02";
      when x"092c" => bus_data_in <= x"e2";
      when x"092d" => bus_data_in <= x"24";
      when x"092e" => bus_data_in <= x"14";
      when x"092f" => bus_data_in <= x"18";
      when x"0930" => bus_data_in <= x"08";
      when x"0934" => bus_data_in <= x"58";
      when x"0935" => bus_data_in <= x"24";
      when x"0936" => bus_data_in <= x"24";
      when x"093a" => bus_data_in <= x"30";
      when x"093b" => bus_data_in <= x"48";
      when x"093c" => bus_data_in <= x"10";
      when x"093d" => bus_data_in <= x"20";
      when x"093e" => bus_data_in <= x"78";
      when x"0944" => bus_data_in <= x"ff";
      when x"0945" => bus_data_in <= x"ff";
      when x"0946" => bus_data_in <= x"ff";
      when x"0947" => bus_data_in <= x"ff";
      when x"0953" => bus_data_in <= x"f3";
      when x"0954" => bus_data_in <= x"31";
      when x"0955" => bus_data_in <= x"ff";
      when x"0956" => bus_data_in <= x"ff";
      when x"0957" => bus_data_in <= x"3e";
      when x"0958" => bus_data_in <= x"e4";
      when x"0959" => bus_data_in <= x"e0";
      when x"095a" => bus_data_in <= x"47";
      when x"095b" => bus_data_in <= x"3e";
      when x"095d" => bus_data_in <= x"e0";
      when x"095e" => bus_data_in <= x"43";
      when x"095f" => bus_data_in <= x"e0";
      when x"0960" => bus_data_in <= x"42";
      when x"0961" => bus_data_in <= x"cd";
      when x"0962" => bus_data_in <= x"9d";
      when x"0963" => bus_data_in <= x"09";
      when x"0964" => bus_data_in <= x"21";
      when x"0965" => bus_data_in <= x"50";
      when x"0966" => bus_data_in <= x"01";
      when x"0967" => bus_data_in <= x"11";
      when x"0969" => bus_data_in <= x"80";
      when x"096a" => bus_data_in <= x"01";
      when x"096c" => bus_data_in <= x"08";
      when x"096d" => bus_data_in <= x"cd";
      when x"096e" => bus_data_in <= x"7b";
      when x"0970" => bus_data_in <= x"3e";
      when x"0971" => bus_data_in <= x"95";
      when x"0972" => bus_data_in <= x"e0";
      when x"0973" => bus_data_in <= x"40";
      when x"0974" => bus_data_in <= x"3e";
      when x"0975" => bus_data_in <= x"20";
      when x"0976" => bus_data_in <= x"21";
      when x"0978" => bus_data_in <= x"98";
      when x"0979" => bus_data_in <= x"01";
      when x"097b" => bus_data_in <= x"04";
      when x"097c" => bus_data_in <= x"cd";
      when x"097d" => bus_data_in <= x"8b";
      when x"097f" => bus_data_in <= x"21";
      when x"0980" => bus_data_in <= x"90";
      when x"0981" => bus_data_in <= x"09";
      when x"0982" => bus_data_in <= x"11";
      when x"0983" => bus_data_in <= x"e3";
      when x"0984" => bus_data_in <= x"98";
      when x"0985" => bus_data_in <= x"01";
      when x"0986" => bus_data_in <= x"0d";
      when x"0988" => bus_data_in <= x"cd";
      when x"0989" => bus_data_in <= x"a1";
      when x"098b" => bus_data_in <= x"76";
      when x"098e" => bus_data_in <= x"18";
      when x"098f" => bus_data_in <= x"fb";
      when x"0990" => bus_data_in <= x"48";
      when x"0991" => bus_data_in <= x"65";
      when x"0992" => bus_data_in <= x"6c";
      when x"0993" => bus_data_in <= x"6c";
      when x"0994" => bus_data_in <= x"6f";
      when x"0995" => bus_data_in <= x"20";
      when x"0996" => bus_data_in <= x"57";
      when x"0997" => bus_data_in <= x"6f";
      when x"0998" => bus_data_in <= x"72";
      when x"0999" => bus_data_in <= x"6c";
      when x"099a" => bus_data_in <= x"64";
      when x"099b" => bus_data_in <= x"20";
      when x"099c" => bus_data_in <= x"21";
      when x"099d" => bus_data_in <= x"f0";
      when x"099e" => bus_data_in <= x"40";
      when x"099f" => bus_data_in <= x"07";
      when x"09a0" => bus_data_in <= x"d0";
      when x"09a1" => bus_data_in <= x"f0";
      when x"09a2" => bus_data_in <= x"44";
      when x"09a3" => bus_data_in <= x"fe";
      when x"09a4" => bus_data_in <= x"91";
      when x"09a5" => bus_data_in <= x"20";
      when x"09a6" => bus_data_in <= x"fa";
      when x"09a7" => bus_data_in <= x"f0";
      when x"09a8" => bus_data_in <= x"40";
      when x"09a9" => bus_data_in <= x"cb";
      when x"09aa" => bus_data_in <= x"bf";
      when x"09ab" => bus_data_in <= x"e0";
      when x"09ac" => bus_data_in <= x"40";
      when x"09ad" => bus_data_in <= x"c9";
      when others => bus_data_in <= x"00";
    end case;
  end process;


  --PREG: process(reset, clock)
  --begin
  --  if reset = '1' then 
  --    ROM_dataout <= x"00";
  --  elsif rising_edge(clock) then 
  --    ROM_dataout <= bus_data_in;
  --  end if;
  --end process;
  --ROM_dataout <= bus_data_in;

  -------------------------------------------------------------------------------
  -- DEVICE UNDER TEST
  -------------------------------------------------------------------------------
  DUT: component processor port map(
    reset => reset,
    clock => clock,

    bus_address => bus_address,
    bus_data_in => bus_data_in,
    bus_data_out => bus_data_out,
    bus_we => bus_we);

  -------------------------------------------------------------------------------
  -- CLOCK
  -------------------------------------------------------------------------------
  PCLK: process
  begin
    clock <= '1';
    wait for clock_period/2;
    clock <= '0';
    wait for clock_period/2;
  end process;
  
end Behavioural;
