library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library work;
use work.PKG_gameboy.ALL;

entity processor_tb is
end processor_tb;

architecture Behavioural of processor_tb is

  signal reset, clock : STD_LOGIC;

  signal ROM_address : STD_LOGIC_VECTOR(15 downto 0);
  signal ROM_dataout_i, ROM_dataout : STD_LOGIC_VECTOR(7 downto 0);

  constant clock_period : time := 250 ns;

begin

  -------------------------------------------------------------------------------
  -- STIMULI
  -------------------------------------------------------------------------------
  PSTIM: process
  begin
    reset <= '1';
    wait for clock_period*2;

    reset <= '0';
    wait for clock_period*2;



    wait;
  end process;

  -------------------------------------------------------------------------------
  -- MEMORY MODEL
  -------------------------------------------------------------------------------
  PMUX: process(ROM_address)
  begin
    case ROM_address is
      when x"0040" => ROM_dataout_i <= x"d9";
      when x"0048" => ROM_dataout_i <= x"d9";
      when x"0050" => ROM_dataout_i <= x"d9";
      when x"0058" => ROM_dataout_i <= x"d9";
      when x"0060" => ROM_dataout_i <= x"d9";
      when x"0061" => ROM_dataout_i <= x"04";
      when x"0062" => ROM_dataout_i <= x"0c";
      when x"0063" => ROM_dataout_i <= x"18";
      when x"0064" => ROM_dataout_i <= x"01";
      when x"0065" => ROM_dataout_i <= x"22";
      when x"0066" => ROM_dataout_i <= x"0d";
      when x"0067" => ROM_dataout_i <= x"20";
      when x"0068" => ROM_dataout_i <= x"fc";
      when x"0069" => ROM_dataout_i <= x"05";
      when x"006a" => ROM_dataout_i <= x"20";
      when x"006b" => ROM_dataout_i <= x"f9";
      when x"006c" => ROM_dataout_i <= x"c9";
      when x"006d" => ROM_dataout_i <= x"04";
      when x"006e" => ROM_dataout_i <= x"0c";
      when x"006f" => ROM_dataout_i <= x"18";
      when x"0070" => ROM_dataout_i <= x"03";
      when x"0071" => ROM_dataout_i <= x"2a";
      when x"0072" => ROM_dataout_i <= x"12";
      when x"0073" => ROM_dataout_i <= x"13";
      when x"0074" => ROM_dataout_i <= x"0d";
      when x"0075" => ROM_dataout_i <= x"20";
      when x"0076" => ROM_dataout_i <= x"fa";
      when x"0077" => ROM_dataout_i <= x"05";
      when x"0078" => ROM_dataout_i <= x"20";
      when x"0079" => ROM_dataout_i <= x"f7";
      when x"007a" => ROM_dataout_i <= x"c9";
      when x"007b" => ROM_dataout_i <= x"04";
      when x"007c" => ROM_dataout_i <= x"0c";
      when x"007d" => ROM_dataout_i <= x"18";
      when x"007e" => ROM_dataout_i <= x"05";
      when x"007f" => ROM_dataout_i <= x"2a";
      when x"0080" => ROM_dataout_i <= x"12";
      when x"0081" => ROM_dataout_i <= x"13";
      when x"0082" => ROM_dataout_i <= x"12";
      when x"0083" => ROM_dataout_i <= x"13";
      when x"0084" => ROM_dataout_i <= x"0d";
      when x"0085" => ROM_dataout_i <= x"20";
      when x"0086" => ROM_dataout_i <= x"f8";
      when x"0087" => ROM_dataout_i <= x"05";
      when x"0088" => ROM_dataout_i <= x"20";
      when x"0089" => ROM_dataout_i <= x"f5";
      when x"008a" => ROM_dataout_i <= x"c9";
      when x"008b" => ROM_dataout_i <= x"04";
      when x"008c" => ROM_dataout_i <= x"0c";
      when x"008d" => ROM_dataout_i <= x"18";
      when x"008e" => ROM_dataout_i <= x"0b";
      when x"008f" => ROM_dataout_i <= x"f5";
      when x"0090" => ROM_dataout_i <= x"f3";
      when x"0091" => ROM_dataout_i <= x"f0";
      when x"0092" => ROM_dataout_i <= x"41";
      when x"0093" => ROM_dataout_i <= x"e6";
      when x"0094" => ROM_dataout_i <= x"02";
      when x"0095" => ROM_dataout_i <= x"20";
      when x"0096" => ROM_dataout_i <= x"fa";
      when x"0097" => ROM_dataout_i <= x"f1";
      when x"0098" => ROM_dataout_i <= x"22";
      when x"0099" => ROM_dataout_i <= x"fb";
      when x"009a" => ROM_dataout_i <= x"0d";
      when x"009b" => ROM_dataout_i <= x"20";
      when x"009c" => ROM_dataout_i <= x"f2";
      when x"009d" => ROM_dataout_i <= x"05";
      when x"009e" => ROM_dataout_i <= x"20";
      when x"009f" => ROM_dataout_i <= x"ef";
      when x"00a0" => ROM_dataout_i <= x"c9";
      when x"00a1" => ROM_dataout_i <= x"04";
      when x"00a2" => ROM_dataout_i <= x"0c";
      when x"00a3" => ROM_dataout_i <= x"18";
      when x"00a4" => ROM_dataout_i <= x"0b";
      when x"00a5" => ROM_dataout_i <= x"f3";
      when x"00a6" => ROM_dataout_i <= x"f0";
      when x"00a7" => ROM_dataout_i <= x"41";
      when x"00a8" => ROM_dataout_i <= x"e6";
      when x"00a9" => ROM_dataout_i <= x"02";
      when x"00aa" => ROM_dataout_i <= x"20";
      when x"00ab" => ROM_dataout_i <= x"fa";
      when x"00ac" => ROM_dataout_i <= x"2a";
      when x"00ad" => ROM_dataout_i <= x"12";
      when x"00ae" => ROM_dataout_i <= x"fb";
      when x"00af" => ROM_dataout_i <= x"13";
      when x"00b0" => ROM_dataout_i <= x"0d";
      when x"00b1" => ROM_dataout_i <= x"20";
      when x"00b2" => ROM_dataout_i <= x"f2";
      when x"00b3" => ROM_dataout_i <= x"05";
      when x"00b4" => ROM_dataout_i <= x"20";
      when x"00b5" => ROM_dataout_i <= x"ef";
      when x"00b6" => ROM_dataout_i <= x"c9";
      when x"0101" => ROM_dataout_i <= x"c3";
      when x"0102" => ROM_dataout_i <= x"52";
      when x"0103" => ROM_dataout_i <= x"09";
      when x"0104" => ROM_dataout_i <= x"ce";
      when x"0105" => ROM_dataout_i <= x"ed";
      when x"0106" => ROM_dataout_i <= x"66";
      when x"0107" => ROM_dataout_i <= x"66";
      when x"0108" => ROM_dataout_i <= x"cc";
      when x"0109" => ROM_dataout_i <= x"0d";
      when x"010b" => ROM_dataout_i <= x"0b";
      when x"010c" => ROM_dataout_i <= x"03";
      when x"010d" => ROM_dataout_i <= x"73";
      when x"010f" => ROM_dataout_i <= x"83";
      when x"0111" => ROM_dataout_i <= x"0c";
      when x"0113" => ROM_dataout_i <= x"0d";
      when x"0115" => ROM_dataout_i <= x"08";
      when x"0116" => ROM_dataout_i <= x"11";
      when x"0117" => ROM_dataout_i <= x"1f";
      when x"0118" => ROM_dataout_i <= x"88";
      when x"0119" => ROM_dataout_i <= x"89";
      when x"011b" => ROM_dataout_i <= x"0e";
      when x"011c" => ROM_dataout_i <= x"dc";
      when x"011d" => ROM_dataout_i <= x"cc";
      when x"011e" => ROM_dataout_i <= x"6e";
      when x"011f" => ROM_dataout_i <= x"e6";
      when x"0120" => ROM_dataout_i <= x"dd";
      when x"0121" => ROM_dataout_i <= x"dd";
      when x"0122" => ROM_dataout_i <= x"d9";
      when x"0123" => ROM_dataout_i <= x"99";
      when x"0124" => ROM_dataout_i <= x"bb";
      when x"0125" => ROM_dataout_i <= x"bb";
      when x"0126" => ROM_dataout_i <= x"67";
      when x"0127" => ROM_dataout_i <= x"63";
      when x"0128" => ROM_dataout_i <= x"6e";
      when x"0129" => ROM_dataout_i <= x"0e";
      when x"012a" => ROM_dataout_i <= x"ec";
      when x"012b" => ROM_dataout_i <= x"cc";
      when x"012c" => ROM_dataout_i <= x"dd";
      when x"012d" => ROM_dataout_i <= x"dc";
      when x"012e" => ROM_dataout_i <= x"99";
      when x"012f" => ROM_dataout_i <= x"9f";
      when x"0130" => ROM_dataout_i <= x"bb";
      when x"0131" => ROM_dataout_i <= x"b9";
      when x"0132" => ROM_dataout_i <= x"33";
      when x"0133" => ROM_dataout_i <= x"3e";
      when x"0134" => ROM_dataout_i <= x"45";
      when x"0135" => ROM_dataout_i <= x"58";
      when x"0136" => ROM_dataout_i <= x"41";
      when x"0137" => ROM_dataout_i <= x"4d";
      when x"0138" => ROM_dataout_i <= x"50";
      when x"0139" => ROM_dataout_i <= x"4c";
      when x"013a" => ROM_dataout_i <= x"45";
      when x"014a" => ROM_dataout_i <= x"01";
      when x"014b" => ROM_dataout_i <= x"33";
      when x"014d" => ROM_dataout_i <= x"a7";
      when x"014e" => ROM_dataout_i <= x"f8";
      when x"014f" => ROM_dataout_i <= x"5f";
      when x"0150" => ROM_dataout_i <= x"7e";
      when x"0151" => ROM_dataout_i <= x"42";
      when x"0152" => ROM_dataout_i <= x"42";
      when x"0153" => ROM_dataout_i <= x"42";
      when x"0154" => ROM_dataout_i <= x"42";
      when x"0155" => ROM_dataout_i <= x"42";
      when x"0156" => ROM_dataout_i <= x"42";
      when x"0157" => ROM_dataout_i <= x"7e";
      when x"0158" => ROM_dataout_i <= x"7e";
      when x"0159" => ROM_dataout_i <= x"81";
      when x"015a" => ROM_dataout_i <= x"a5";
      when x"015b" => ROM_dataout_i <= x"81";
      when x"015c" => ROM_dataout_i <= x"bd";
      when x"015d" => ROM_dataout_i <= x"99";
      when x"015e" => ROM_dataout_i <= x"81";
      when x"015f" => ROM_dataout_i <= x"7e";
      when x"0160" => ROM_dataout_i <= x"7e";
      when x"0161" => ROM_dataout_i <= x"ff";
      when x"0162" => ROM_dataout_i <= x"db";
      when x"0163" => ROM_dataout_i <= x"ff";
      when x"0164" => ROM_dataout_i <= x"c3";
      when x"0165" => ROM_dataout_i <= x"e7";
      when x"0166" => ROM_dataout_i <= x"ff";
      when x"0167" => ROM_dataout_i <= x"7e";
      when x"0168" => ROM_dataout_i <= x"6c";
      when x"0169" => ROM_dataout_i <= x"fe";
      when x"016a" => ROM_dataout_i <= x"fe";
      when x"016b" => ROM_dataout_i <= x"fe";
      when x"016c" => ROM_dataout_i <= x"7c";
      when x"016d" => ROM_dataout_i <= x"38";
      when x"016e" => ROM_dataout_i <= x"10";
      when x"0170" => ROM_dataout_i <= x"10";
      when x"0171" => ROM_dataout_i <= x"38";
      when x"0172" => ROM_dataout_i <= x"7c";
      when x"0173" => ROM_dataout_i <= x"fe";
      when x"0174" => ROM_dataout_i <= x"7c";
      when x"0175" => ROM_dataout_i <= x"38";
      when x"0176" => ROM_dataout_i <= x"10";
      when x"0178" => ROM_dataout_i <= x"38";
      when x"0179" => ROM_dataout_i <= x"7c";
      when x"017a" => ROM_dataout_i <= x"38";
      when x"017b" => ROM_dataout_i <= x"fe";
      when x"017c" => ROM_dataout_i <= x"fe";
      when x"017d" => ROM_dataout_i <= x"7c";
      when x"017e" => ROM_dataout_i <= x"38";
      when x"017f" => ROM_dataout_i <= x"7c";
      when x"0180" => ROM_dataout_i <= x"10";
      when x"0181" => ROM_dataout_i <= x"10";
      when x"0182" => ROM_dataout_i <= x"38";
      when x"0183" => ROM_dataout_i <= x"7c";
      when x"0184" => ROM_dataout_i <= x"fe";
      when x"0185" => ROM_dataout_i <= x"7c";
      when x"0186" => ROM_dataout_i <= x"38";
      when x"0187" => ROM_dataout_i <= x"7c";
      when x"018a" => ROM_dataout_i <= x"18";
      when x"018b" => ROM_dataout_i <= x"3c";
      when x"018c" => ROM_dataout_i <= x"3c";
      when x"018d" => ROM_dataout_i <= x"18";
      when x"0190" => ROM_dataout_i <= x"ff";
      when x"0191" => ROM_dataout_i <= x"ff";
      when x"0192" => ROM_dataout_i <= x"e7";
      when x"0193" => ROM_dataout_i <= x"c3";
      when x"0194" => ROM_dataout_i <= x"c3";
      when x"0195" => ROM_dataout_i <= x"e7";
      when x"0196" => ROM_dataout_i <= x"ff";
      when x"0197" => ROM_dataout_i <= x"ff";
      when x"0199" => ROM_dataout_i <= x"3c";
      when x"019a" => ROM_dataout_i <= x"66";
      when x"019b" => ROM_dataout_i <= x"42";
      when x"019c" => ROM_dataout_i <= x"42";
      when x"019d" => ROM_dataout_i <= x"66";
      when x"019e" => ROM_dataout_i <= x"3c";
      when x"01a0" => ROM_dataout_i <= x"ff";
      when x"01a1" => ROM_dataout_i <= x"c3";
      when x"01a2" => ROM_dataout_i <= x"99";
      when x"01a3" => ROM_dataout_i <= x"bd";
      when x"01a4" => ROM_dataout_i <= x"bd";
      when x"01a5" => ROM_dataout_i <= x"99";
      when x"01a6" => ROM_dataout_i <= x"c3";
      when x"01a7" => ROM_dataout_i <= x"ff";
      when x"01a8" => ROM_dataout_i <= x"0f";
      when x"01a9" => ROM_dataout_i <= x"07";
      when x"01aa" => ROM_dataout_i <= x"0f";
      when x"01ab" => ROM_dataout_i <= x"7d";
      when x"01ac" => ROM_dataout_i <= x"cc";
      when x"01ad" => ROM_dataout_i <= x"cc";
      when x"01ae" => ROM_dataout_i <= x"cc";
      when x"01af" => ROM_dataout_i <= x"78";
      when x"01b0" => ROM_dataout_i <= x"3c";
      when x"01b1" => ROM_dataout_i <= x"66";
      when x"01b2" => ROM_dataout_i <= x"66";
      when x"01b3" => ROM_dataout_i <= x"66";
      when x"01b4" => ROM_dataout_i <= x"3c";
      when x"01b5" => ROM_dataout_i <= x"18";
      when x"01b6" => ROM_dataout_i <= x"7e";
      when x"01b7" => ROM_dataout_i <= x"18";
      when x"01b8" => ROM_dataout_i <= x"3f";
      when x"01b9" => ROM_dataout_i <= x"33";
      when x"01ba" => ROM_dataout_i <= x"3f";
      when x"01bb" => ROM_dataout_i <= x"30";
      when x"01bc" => ROM_dataout_i <= x"30";
      when x"01bd" => ROM_dataout_i <= x"70";
      when x"01be" => ROM_dataout_i <= x"f0";
      when x"01bf" => ROM_dataout_i <= x"e0";
      when x"01c0" => ROM_dataout_i <= x"7f";
      when x"01c1" => ROM_dataout_i <= x"63";
      when x"01c2" => ROM_dataout_i <= x"7f";
      when x"01c3" => ROM_dataout_i <= x"63";
      when x"01c4" => ROM_dataout_i <= x"63";
      when x"01c5" => ROM_dataout_i <= x"67";
      when x"01c6" => ROM_dataout_i <= x"e6";
      when x"01c7" => ROM_dataout_i <= x"c0";
      when x"01c8" => ROM_dataout_i <= x"99";
      when x"01c9" => ROM_dataout_i <= x"5a";
      when x"01ca" => ROM_dataout_i <= x"3c";
      when x"01cb" => ROM_dataout_i <= x"e7";
      when x"01cc" => ROM_dataout_i <= x"e7";
      when x"01cd" => ROM_dataout_i <= x"3c";
      when x"01ce" => ROM_dataout_i <= x"5a";
      when x"01cf" => ROM_dataout_i <= x"99";
      when x"01d0" => ROM_dataout_i <= x"80";
      when x"01d1" => ROM_dataout_i <= x"e0";
      when x"01d2" => ROM_dataout_i <= x"f8";
      when x"01d3" => ROM_dataout_i <= x"fe";
      when x"01d4" => ROM_dataout_i <= x"f8";
      when x"01d5" => ROM_dataout_i <= x"e0";
      when x"01d6" => ROM_dataout_i <= x"80";
      when x"01d8" => ROM_dataout_i <= x"02";
      when x"01d9" => ROM_dataout_i <= x"0e";
      when x"01da" => ROM_dataout_i <= x"3e";
      when x"01db" => ROM_dataout_i <= x"fe";
      when x"01dc" => ROM_dataout_i <= x"3e";
      when x"01dd" => ROM_dataout_i <= x"0e";
      when x"01de" => ROM_dataout_i <= x"02";
      when x"01e0" => ROM_dataout_i <= x"18";
      when x"01e1" => ROM_dataout_i <= x"3c";
      when x"01e2" => ROM_dataout_i <= x"7e";
      when x"01e3" => ROM_dataout_i <= x"18";
      when x"01e4" => ROM_dataout_i <= x"18";
      when x"01e5" => ROM_dataout_i <= x"7e";
      when x"01e6" => ROM_dataout_i <= x"3c";
      when x"01e7" => ROM_dataout_i <= x"18";
      when x"01e8" => ROM_dataout_i <= x"66";
      when x"01e9" => ROM_dataout_i <= x"66";
      when x"01ea" => ROM_dataout_i <= x"66";
      when x"01eb" => ROM_dataout_i <= x"66";
      when x"01ec" => ROM_dataout_i <= x"66";
      when x"01ee" => ROM_dataout_i <= x"66";
      when x"01f0" => ROM_dataout_i <= x"7f";
      when x"01f1" => ROM_dataout_i <= x"db";
      when x"01f2" => ROM_dataout_i <= x"db";
      when x"01f3" => ROM_dataout_i <= x"7b";
      when x"01f4" => ROM_dataout_i <= x"1b";
      when x"01f5" => ROM_dataout_i <= x"1b";
      when x"01f6" => ROM_dataout_i <= x"1b";
      when x"01f8" => ROM_dataout_i <= x"3e";
      when x"01f9" => ROM_dataout_i <= x"63";
      when x"01fa" => ROM_dataout_i <= x"38";
      when x"01fb" => ROM_dataout_i <= x"6c";
      when x"01fc" => ROM_dataout_i <= x"6c";
      when x"01fd" => ROM_dataout_i <= x"38";
      when x"01fe" => ROM_dataout_i <= x"cc";
      when x"01ff" => ROM_dataout_i <= x"78";
      when x"0204" => ROM_dataout_i <= x"7e";
      when x"0205" => ROM_dataout_i <= x"7e";
      when x"0206" => ROM_dataout_i <= x"7e";
      when x"0208" => ROM_dataout_i <= x"18";
      when x"0209" => ROM_dataout_i <= x"3c";
      when x"020a" => ROM_dataout_i <= x"7e";
      when x"020b" => ROM_dataout_i <= x"18";
      when x"020c" => ROM_dataout_i <= x"7e";
      when x"020d" => ROM_dataout_i <= x"3c";
      when x"020e" => ROM_dataout_i <= x"18";
      when x"020f" => ROM_dataout_i <= x"ff";
      when x"0210" => ROM_dataout_i <= x"18";
      when x"0211" => ROM_dataout_i <= x"3c";
      when x"0212" => ROM_dataout_i <= x"7e";
      when x"0213" => ROM_dataout_i <= x"18";
      when x"0214" => ROM_dataout_i <= x"18";
      when x"0215" => ROM_dataout_i <= x"18";
      when x"0216" => ROM_dataout_i <= x"18";
      when x"0218" => ROM_dataout_i <= x"18";
      when x"0219" => ROM_dataout_i <= x"18";
      when x"021a" => ROM_dataout_i <= x"18";
      when x"021b" => ROM_dataout_i <= x"18";
      when x"021c" => ROM_dataout_i <= x"7e";
      when x"021d" => ROM_dataout_i <= x"3c";
      when x"021e" => ROM_dataout_i <= x"18";
      when x"0221" => ROM_dataout_i <= x"18";
      when x"0222" => ROM_dataout_i <= x"0c";
      when x"0223" => ROM_dataout_i <= x"fe";
      when x"0224" => ROM_dataout_i <= x"0c";
      when x"0225" => ROM_dataout_i <= x"18";
      when x"0229" => ROM_dataout_i <= x"30";
      when x"022a" => ROM_dataout_i <= x"60";
      when x"022b" => ROM_dataout_i <= x"fe";
      when x"022c" => ROM_dataout_i <= x"60";
      when x"022d" => ROM_dataout_i <= x"30";
      when x"0232" => ROM_dataout_i <= x"c0";
      when x"0233" => ROM_dataout_i <= x"c0";
      when x"0234" => ROM_dataout_i <= x"c0";
      when x"0235" => ROM_dataout_i <= x"fe";
      when x"0239" => ROM_dataout_i <= x"24";
      when x"023a" => ROM_dataout_i <= x"66";
      when x"023b" => ROM_dataout_i <= x"ff";
      when x"023c" => ROM_dataout_i <= x"66";
      when x"023d" => ROM_dataout_i <= x"24";
      when x"0241" => ROM_dataout_i <= x"18";
      when x"0242" => ROM_dataout_i <= x"3c";
      when x"0243" => ROM_dataout_i <= x"7e";
      when x"0244" => ROM_dataout_i <= x"ff";
      when x"0245" => ROM_dataout_i <= x"ff";
      when x"0249" => ROM_dataout_i <= x"ff";
      when x"024a" => ROM_dataout_i <= x"ff";
      when x"024b" => ROM_dataout_i <= x"7e";
      when x"024c" => ROM_dataout_i <= x"3c";
      when x"024d" => ROM_dataout_i <= x"18";
      when x"0258" => ROM_dataout_i <= x"30";
      when x"0259" => ROM_dataout_i <= x"30";
      when x"025a" => ROM_dataout_i <= x"30";
      when x"025b" => ROM_dataout_i <= x"30";
      when x"025c" => ROM_dataout_i <= x"30";
      when x"025e" => ROM_dataout_i <= x"30";
      when x"0260" => ROM_dataout_i <= x"6c";
      when x"0261" => ROM_dataout_i <= x"6c";
      when x"0262" => ROM_dataout_i <= x"6c";
      when x"0268" => ROM_dataout_i <= x"6c";
      when x"0269" => ROM_dataout_i <= x"6c";
      when x"026a" => ROM_dataout_i <= x"fe";
      when x"026b" => ROM_dataout_i <= x"6c";
      when x"026c" => ROM_dataout_i <= x"fe";
      when x"026d" => ROM_dataout_i <= x"6c";
      when x"026e" => ROM_dataout_i <= x"6c";
      when x"0270" => ROM_dataout_i <= x"30";
      when x"0271" => ROM_dataout_i <= x"7c";
      when x"0272" => ROM_dataout_i <= x"c0";
      when x"0273" => ROM_dataout_i <= x"78";
      when x"0274" => ROM_dataout_i <= x"0c";
      when x"0275" => ROM_dataout_i <= x"f8";
      when x"0276" => ROM_dataout_i <= x"30";
      when x"0279" => ROM_dataout_i <= x"c6";
      when x"027a" => ROM_dataout_i <= x"cc";
      when x"027b" => ROM_dataout_i <= x"18";
      when x"027c" => ROM_dataout_i <= x"30";
      when x"027d" => ROM_dataout_i <= x"66";
      when x"027e" => ROM_dataout_i <= x"c6";
      when x"0280" => ROM_dataout_i <= x"38";
      when x"0281" => ROM_dataout_i <= x"6c";
      when x"0282" => ROM_dataout_i <= x"38";
      when x"0283" => ROM_dataout_i <= x"76";
      when x"0284" => ROM_dataout_i <= x"dc";
      when x"0285" => ROM_dataout_i <= x"cc";
      when x"0286" => ROM_dataout_i <= x"76";
      when x"0288" => ROM_dataout_i <= x"60";
      when x"0289" => ROM_dataout_i <= x"60";
      when x"028a" => ROM_dataout_i <= x"c0";
      when x"0290" => ROM_dataout_i <= x"18";
      when x"0291" => ROM_dataout_i <= x"30";
      when x"0292" => ROM_dataout_i <= x"60";
      when x"0293" => ROM_dataout_i <= x"60";
      when x"0294" => ROM_dataout_i <= x"60";
      when x"0295" => ROM_dataout_i <= x"30";
      when x"0296" => ROM_dataout_i <= x"18";
      when x"0298" => ROM_dataout_i <= x"60";
      when x"0299" => ROM_dataout_i <= x"30";
      when x"029a" => ROM_dataout_i <= x"18";
      when x"029b" => ROM_dataout_i <= x"18";
      when x"029c" => ROM_dataout_i <= x"18";
      when x"029d" => ROM_dataout_i <= x"30";
      when x"029e" => ROM_dataout_i <= x"60";
      when x"02a1" => ROM_dataout_i <= x"66";
      when x"02a2" => ROM_dataout_i <= x"3c";
      when x"02a3" => ROM_dataout_i <= x"ff";
      when x"02a4" => ROM_dataout_i <= x"3c";
      when x"02a5" => ROM_dataout_i <= x"66";
      when x"02a9" => ROM_dataout_i <= x"30";
      when x"02aa" => ROM_dataout_i <= x"30";
      when x"02ab" => ROM_dataout_i <= x"fc";
      when x"02ac" => ROM_dataout_i <= x"30";
      when x"02ad" => ROM_dataout_i <= x"30";
      when x"02b5" => ROM_dataout_i <= x"30";
      when x"02b6" => ROM_dataout_i <= x"30";
      when x"02b7" => ROM_dataout_i <= x"60";
      when x"02bb" => ROM_dataout_i <= x"fc";
      when x"02c5" => ROM_dataout_i <= x"30";
      when x"02c6" => ROM_dataout_i <= x"30";
      when x"02c8" => ROM_dataout_i <= x"06";
      when x"02c9" => ROM_dataout_i <= x"0c";
      when x"02ca" => ROM_dataout_i <= x"18";
      when x"02cb" => ROM_dataout_i <= x"30";
      when x"02cc" => ROM_dataout_i <= x"60";
      when x"02cd" => ROM_dataout_i <= x"c0";
      when x"02ce" => ROM_dataout_i <= x"80";
      when x"02d0" => ROM_dataout_i <= x"7c";
      when x"02d1" => ROM_dataout_i <= x"c6";
      when x"02d2" => ROM_dataout_i <= x"ce";
      when x"02d3" => ROM_dataout_i <= x"de";
      when x"02d4" => ROM_dataout_i <= x"f6";
      when x"02d5" => ROM_dataout_i <= x"e6";
      when x"02d6" => ROM_dataout_i <= x"7c";
      when x"02d8" => ROM_dataout_i <= x"30";
      when x"02d9" => ROM_dataout_i <= x"70";
      when x"02da" => ROM_dataout_i <= x"30";
      when x"02db" => ROM_dataout_i <= x"30";
      when x"02dc" => ROM_dataout_i <= x"30";
      when x"02dd" => ROM_dataout_i <= x"30";
      when x"02de" => ROM_dataout_i <= x"fc";
      when x"02e0" => ROM_dataout_i <= x"78";
      when x"02e1" => ROM_dataout_i <= x"cc";
      when x"02e2" => ROM_dataout_i <= x"0c";
      when x"02e3" => ROM_dataout_i <= x"38";
      when x"02e4" => ROM_dataout_i <= x"60";
      when x"02e5" => ROM_dataout_i <= x"cc";
      when x"02e6" => ROM_dataout_i <= x"fc";
      when x"02e8" => ROM_dataout_i <= x"78";
      when x"02e9" => ROM_dataout_i <= x"cc";
      when x"02ea" => ROM_dataout_i <= x"0c";
      when x"02eb" => ROM_dataout_i <= x"38";
      when x"02ec" => ROM_dataout_i <= x"0c";
      when x"02ed" => ROM_dataout_i <= x"cc";
      when x"02ee" => ROM_dataout_i <= x"78";
      when x"02f0" => ROM_dataout_i <= x"1c";
      when x"02f1" => ROM_dataout_i <= x"3c";
      when x"02f2" => ROM_dataout_i <= x"6c";
      when x"02f3" => ROM_dataout_i <= x"cc";
      when x"02f4" => ROM_dataout_i <= x"fe";
      when x"02f5" => ROM_dataout_i <= x"0c";
      when x"02f6" => ROM_dataout_i <= x"1e";
      when x"02f8" => ROM_dataout_i <= x"fc";
      when x"02f9" => ROM_dataout_i <= x"c0";
      when x"02fa" => ROM_dataout_i <= x"f8";
      when x"02fb" => ROM_dataout_i <= x"0c";
      when x"02fc" => ROM_dataout_i <= x"0c";
      when x"02fd" => ROM_dataout_i <= x"cc";
      when x"02fe" => ROM_dataout_i <= x"78";
      when x"0300" => ROM_dataout_i <= x"38";
      when x"0301" => ROM_dataout_i <= x"60";
      when x"0302" => ROM_dataout_i <= x"c0";
      when x"0303" => ROM_dataout_i <= x"f8";
      when x"0304" => ROM_dataout_i <= x"cc";
      when x"0305" => ROM_dataout_i <= x"cc";
      when x"0306" => ROM_dataout_i <= x"78";
      when x"0308" => ROM_dataout_i <= x"fc";
      when x"0309" => ROM_dataout_i <= x"cc";
      when x"030a" => ROM_dataout_i <= x"0c";
      when x"030b" => ROM_dataout_i <= x"18";
      when x"030c" => ROM_dataout_i <= x"30";
      when x"030d" => ROM_dataout_i <= x"30";
      when x"030e" => ROM_dataout_i <= x"30";
      when x"0310" => ROM_dataout_i <= x"78";
      when x"0311" => ROM_dataout_i <= x"cc";
      when x"0312" => ROM_dataout_i <= x"cc";
      when x"0313" => ROM_dataout_i <= x"78";
      when x"0314" => ROM_dataout_i <= x"cc";
      when x"0315" => ROM_dataout_i <= x"cc";
      when x"0316" => ROM_dataout_i <= x"78";
      when x"0318" => ROM_dataout_i <= x"78";
      when x"0319" => ROM_dataout_i <= x"cc";
      when x"031a" => ROM_dataout_i <= x"cc";
      when x"031b" => ROM_dataout_i <= x"7c";
      when x"031c" => ROM_dataout_i <= x"0c";
      when x"031d" => ROM_dataout_i <= x"18";
      when x"031e" => ROM_dataout_i <= x"70";
      when x"0321" => ROM_dataout_i <= x"30";
      when x"0322" => ROM_dataout_i <= x"30";
      when x"0325" => ROM_dataout_i <= x"30";
      when x"0326" => ROM_dataout_i <= x"30";
      when x"0329" => ROM_dataout_i <= x"30";
      when x"032a" => ROM_dataout_i <= x"30";
      when x"032d" => ROM_dataout_i <= x"30";
      when x"032e" => ROM_dataout_i <= x"30";
      when x"032f" => ROM_dataout_i <= x"60";
      when x"0330" => ROM_dataout_i <= x"18";
      when x"0331" => ROM_dataout_i <= x"30";
      when x"0332" => ROM_dataout_i <= x"60";
      when x"0333" => ROM_dataout_i <= x"c0";
      when x"0334" => ROM_dataout_i <= x"60";
      when x"0335" => ROM_dataout_i <= x"30";
      when x"0336" => ROM_dataout_i <= x"18";
      when x"033a" => ROM_dataout_i <= x"fc";
      when x"033d" => ROM_dataout_i <= x"fc";
      when x"0340" => ROM_dataout_i <= x"60";
      when x"0341" => ROM_dataout_i <= x"30";
      when x"0342" => ROM_dataout_i <= x"18";
      when x"0343" => ROM_dataout_i <= x"0c";
      when x"0344" => ROM_dataout_i <= x"18";
      when x"0345" => ROM_dataout_i <= x"30";
      when x"0346" => ROM_dataout_i <= x"60";
      when x"0348" => ROM_dataout_i <= x"78";
      when x"0349" => ROM_dataout_i <= x"cc";
      when x"034a" => ROM_dataout_i <= x"0c";
      when x"034b" => ROM_dataout_i <= x"18";
      when x"034c" => ROM_dataout_i <= x"30";
      when x"034e" => ROM_dataout_i <= x"30";
      when x"0350" => ROM_dataout_i <= x"7c";
      when x"0351" => ROM_dataout_i <= x"c6";
      when x"0352" => ROM_dataout_i <= x"de";
      when x"0353" => ROM_dataout_i <= x"de";
      when x"0354" => ROM_dataout_i <= x"de";
      when x"0355" => ROM_dataout_i <= x"c0";
      when x"0356" => ROM_dataout_i <= x"78";
      when x"0358" => ROM_dataout_i <= x"30";
      when x"0359" => ROM_dataout_i <= x"78";
      when x"035a" => ROM_dataout_i <= x"cc";
      when x"035b" => ROM_dataout_i <= x"cc";
      when x"035c" => ROM_dataout_i <= x"fc";
      when x"035d" => ROM_dataout_i <= x"cc";
      when x"035e" => ROM_dataout_i <= x"cc";
      when x"0360" => ROM_dataout_i <= x"fc";
      when x"0361" => ROM_dataout_i <= x"66";
      when x"0362" => ROM_dataout_i <= x"66";
      when x"0363" => ROM_dataout_i <= x"7c";
      when x"0364" => ROM_dataout_i <= x"66";
      when x"0365" => ROM_dataout_i <= x"66";
      when x"0366" => ROM_dataout_i <= x"fc";
      when x"0368" => ROM_dataout_i <= x"3c";
      when x"0369" => ROM_dataout_i <= x"66";
      when x"036a" => ROM_dataout_i <= x"c0";
      when x"036b" => ROM_dataout_i <= x"c0";
      when x"036c" => ROM_dataout_i <= x"c0";
      when x"036d" => ROM_dataout_i <= x"66";
      when x"036e" => ROM_dataout_i <= x"3c";
      when x"0370" => ROM_dataout_i <= x"f8";
      when x"0371" => ROM_dataout_i <= x"6c";
      when x"0372" => ROM_dataout_i <= x"66";
      when x"0373" => ROM_dataout_i <= x"66";
      when x"0374" => ROM_dataout_i <= x"66";
      when x"0375" => ROM_dataout_i <= x"6c";
      when x"0376" => ROM_dataout_i <= x"f8";
      when x"0378" => ROM_dataout_i <= x"7e";
      when x"0379" => ROM_dataout_i <= x"60";
      when x"037a" => ROM_dataout_i <= x"60";
      when x"037b" => ROM_dataout_i <= x"78";
      when x"037c" => ROM_dataout_i <= x"60";
      when x"037d" => ROM_dataout_i <= x"60";
      when x"037e" => ROM_dataout_i <= x"7e";
      when x"0380" => ROM_dataout_i <= x"7e";
      when x"0381" => ROM_dataout_i <= x"60";
      when x"0382" => ROM_dataout_i <= x"60";
      when x"0383" => ROM_dataout_i <= x"78";
      when x"0384" => ROM_dataout_i <= x"60";
      when x"0385" => ROM_dataout_i <= x"60";
      when x"0386" => ROM_dataout_i <= x"60";
      when x"0388" => ROM_dataout_i <= x"3c";
      when x"0389" => ROM_dataout_i <= x"66";
      when x"038a" => ROM_dataout_i <= x"c0";
      when x"038b" => ROM_dataout_i <= x"c0";
      when x"038c" => ROM_dataout_i <= x"ce";
      when x"038d" => ROM_dataout_i <= x"66";
      when x"038e" => ROM_dataout_i <= x"3e";
      when x"0390" => ROM_dataout_i <= x"cc";
      when x"0391" => ROM_dataout_i <= x"cc";
      when x"0392" => ROM_dataout_i <= x"cc";
      when x"0393" => ROM_dataout_i <= x"fc";
      when x"0394" => ROM_dataout_i <= x"cc";
      when x"0395" => ROM_dataout_i <= x"cc";
      when x"0396" => ROM_dataout_i <= x"cc";
      when x"0398" => ROM_dataout_i <= x"78";
      when x"0399" => ROM_dataout_i <= x"30";
      when x"039a" => ROM_dataout_i <= x"30";
      when x"039b" => ROM_dataout_i <= x"30";
      when x"039c" => ROM_dataout_i <= x"30";
      when x"039d" => ROM_dataout_i <= x"30";
      when x"039e" => ROM_dataout_i <= x"78";
      when x"03a0" => ROM_dataout_i <= x"1e";
      when x"03a1" => ROM_dataout_i <= x"0c";
      when x"03a2" => ROM_dataout_i <= x"0c";
      when x"03a3" => ROM_dataout_i <= x"0c";
      when x"03a4" => ROM_dataout_i <= x"cc";
      when x"03a5" => ROM_dataout_i <= x"cc";
      when x"03a6" => ROM_dataout_i <= x"78";
      when x"03a8" => ROM_dataout_i <= x"e6";
      when x"03a9" => ROM_dataout_i <= x"66";
      when x"03aa" => ROM_dataout_i <= x"6c";
      when x"03ab" => ROM_dataout_i <= x"78";
      when x"03ac" => ROM_dataout_i <= x"6c";
      when x"03ad" => ROM_dataout_i <= x"66";
      when x"03ae" => ROM_dataout_i <= x"e6";
      when x"03b0" => ROM_dataout_i <= x"60";
      when x"03b1" => ROM_dataout_i <= x"60";
      when x"03b2" => ROM_dataout_i <= x"60";
      when x"03b3" => ROM_dataout_i <= x"60";
      when x"03b4" => ROM_dataout_i <= x"60";
      when x"03b5" => ROM_dataout_i <= x"60";
      when x"03b6" => ROM_dataout_i <= x"7e";
      when x"03b8" => ROM_dataout_i <= x"c6";
      when x"03b9" => ROM_dataout_i <= x"ee";
      when x"03ba" => ROM_dataout_i <= x"fe";
      when x"03bb" => ROM_dataout_i <= x"fe";
      when x"03bc" => ROM_dataout_i <= x"d6";
      when x"03bd" => ROM_dataout_i <= x"c6";
      when x"03be" => ROM_dataout_i <= x"c6";
      when x"03c0" => ROM_dataout_i <= x"c6";
      when x"03c1" => ROM_dataout_i <= x"e6";
      when x"03c2" => ROM_dataout_i <= x"f6";
      when x"03c3" => ROM_dataout_i <= x"de";
      when x"03c4" => ROM_dataout_i <= x"ce";
      when x"03c5" => ROM_dataout_i <= x"c6";
      when x"03c6" => ROM_dataout_i <= x"c6";
      when x"03c8" => ROM_dataout_i <= x"38";
      when x"03c9" => ROM_dataout_i <= x"6c";
      when x"03ca" => ROM_dataout_i <= x"c6";
      when x"03cb" => ROM_dataout_i <= x"c6";
      when x"03cc" => ROM_dataout_i <= x"c6";
      when x"03cd" => ROM_dataout_i <= x"6c";
      when x"03ce" => ROM_dataout_i <= x"38";
      when x"03d0" => ROM_dataout_i <= x"fc";
      when x"03d1" => ROM_dataout_i <= x"66";
      when x"03d2" => ROM_dataout_i <= x"66";
      when x"03d3" => ROM_dataout_i <= x"7c";
      when x"03d4" => ROM_dataout_i <= x"60";
      when x"03d5" => ROM_dataout_i <= x"60";
      when x"03d6" => ROM_dataout_i <= x"f0";
      when x"03d8" => ROM_dataout_i <= x"78";
      when x"03d9" => ROM_dataout_i <= x"cc";
      when x"03da" => ROM_dataout_i <= x"cc";
      when x"03db" => ROM_dataout_i <= x"cc";
      when x"03dc" => ROM_dataout_i <= x"dc";
      when x"03dd" => ROM_dataout_i <= x"78";
      when x"03de" => ROM_dataout_i <= x"1c";
      when x"03e0" => ROM_dataout_i <= x"fc";
      when x"03e1" => ROM_dataout_i <= x"66";
      when x"03e2" => ROM_dataout_i <= x"66";
      when x"03e3" => ROM_dataout_i <= x"7c";
      when x"03e4" => ROM_dataout_i <= x"6c";
      when x"03e5" => ROM_dataout_i <= x"66";
      when x"03e6" => ROM_dataout_i <= x"e6";
      when x"03e8" => ROM_dataout_i <= x"78";
      when x"03e9" => ROM_dataout_i <= x"cc";
      when x"03ea" => ROM_dataout_i <= x"e0";
      when x"03eb" => ROM_dataout_i <= x"78";
      when x"03ec" => ROM_dataout_i <= x"1c";
      when x"03ed" => ROM_dataout_i <= x"cc";
      when x"03ee" => ROM_dataout_i <= x"78";
      when x"03f0" => ROM_dataout_i <= x"fc";
      when x"03f1" => ROM_dataout_i <= x"30";
      when x"03f2" => ROM_dataout_i <= x"30";
      when x"03f3" => ROM_dataout_i <= x"30";
      when x"03f4" => ROM_dataout_i <= x"30";
      when x"03f5" => ROM_dataout_i <= x"30";
      when x"03f6" => ROM_dataout_i <= x"30";
      when x"03f8" => ROM_dataout_i <= x"cc";
      when x"03f9" => ROM_dataout_i <= x"cc";
      when x"03fa" => ROM_dataout_i <= x"cc";
      when x"03fb" => ROM_dataout_i <= x"cc";
      when x"03fc" => ROM_dataout_i <= x"cc";
      when x"03fd" => ROM_dataout_i <= x"cc";
      when x"03fe" => ROM_dataout_i <= x"fc";
      when x"0400" => ROM_dataout_i <= x"cc";
      when x"0401" => ROM_dataout_i <= x"cc";
      when x"0402" => ROM_dataout_i <= x"cc";
      when x"0403" => ROM_dataout_i <= x"cc";
      when x"0404" => ROM_dataout_i <= x"cc";
      when x"0405" => ROM_dataout_i <= x"78";
      when x"0406" => ROM_dataout_i <= x"30";
      when x"0408" => ROM_dataout_i <= x"c6";
      when x"0409" => ROM_dataout_i <= x"c6";
      when x"040a" => ROM_dataout_i <= x"c6";
      when x"040b" => ROM_dataout_i <= x"d6";
      when x"040c" => ROM_dataout_i <= x"fe";
      when x"040d" => ROM_dataout_i <= x"ee";
      when x"040e" => ROM_dataout_i <= x"c6";
      when x"0410" => ROM_dataout_i <= x"c6";
      when x"0411" => ROM_dataout_i <= x"c6";
      when x"0412" => ROM_dataout_i <= x"6c";
      when x"0413" => ROM_dataout_i <= x"38";
      when x"0414" => ROM_dataout_i <= x"38";
      when x"0415" => ROM_dataout_i <= x"6c";
      when x"0416" => ROM_dataout_i <= x"c6";
      when x"0418" => ROM_dataout_i <= x"cc";
      when x"0419" => ROM_dataout_i <= x"cc";
      when x"041a" => ROM_dataout_i <= x"cc";
      when x"041b" => ROM_dataout_i <= x"78";
      when x"041c" => ROM_dataout_i <= x"30";
      when x"041d" => ROM_dataout_i <= x"30";
      when x"041e" => ROM_dataout_i <= x"78";
      when x"0420" => ROM_dataout_i <= x"fe";
      when x"0421" => ROM_dataout_i <= x"06";
      when x"0422" => ROM_dataout_i <= x"0c";
      when x"0423" => ROM_dataout_i <= x"18";
      when x"0424" => ROM_dataout_i <= x"30";
      when x"0425" => ROM_dataout_i <= x"60";
      when x"0426" => ROM_dataout_i <= x"fe";
      when x"0428" => ROM_dataout_i <= x"78";
      when x"0429" => ROM_dataout_i <= x"60";
      when x"042a" => ROM_dataout_i <= x"60";
      when x"042b" => ROM_dataout_i <= x"60";
      when x"042c" => ROM_dataout_i <= x"60";
      when x"042d" => ROM_dataout_i <= x"60";
      when x"042e" => ROM_dataout_i <= x"78";
      when x"0430" => ROM_dataout_i <= x"c0";
      when x"0431" => ROM_dataout_i <= x"60";
      when x"0432" => ROM_dataout_i <= x"30";
      when x"0433" => ROM_dataout_i <= x"18";
      when x"0434" => ROM_dataout_i <= x"0c";
      when x"0435" => ROM_dataout_i <= x"06";
      when x"0436" => ROM_dataout_i <= x"02";
      when x"0438" => ROM_dataout_i <= x"78";
      when x"0439" => ROM_dataout_i <= x"18";
      when x"043a" => ROM_dataout_i <= x"18";
      when x"043b" => ROM_dataout_i <= x"18";
      when x"043c" => ROM_dataout_i <= x"18";
      when x"043d" => ROM_dataout_i <= x"18";
      when x"043e" => ROM_dataout_i <= x"78";
      when x"0440" => ROM_dataout_i <= x"10";
      when x"0441" => ROM_dataout_i <= x"38";
      when x"0442" => ROM_dataout_i <= x"6c";
      when x"0443" => ROM_dataout_i <= x"c6";
      when x"044f" => ROM_dataout_i <= x"ff";
      when x"0450" => ROM_dataout_i <= x"30";
      when x"0451" => ROM_dataout_i <= x"30";
      when x"0452" => ROM_dataout_i <= x"18";
      when x"045a" => ROM_dataout_i <= x"78";
      when x"045b" => ROM_dataout_i <= x"0c";
      when x"045c" => ROM_dataout_i <= x"7c";
      when x"045d" => ROM_dataout_i <= x"cc";
      when x"045e" => ROM_dataout_i <= x"76";
      when x"0460" => ROM_dataout_i <= x"e0";
      when x"0461" => ROM_dataout_i <= x"60";
      when x"0462" => ROM_dataout_i <= x"60";
      when x"0463" => ROM_dataout_i <= x"7c";
      when x"0464" => ROM_dataout_i <= x"66";
      when x"0465" => ROM_dataout_i <= x"66";
      when x"0466" => ROM_dataout_i <= x"dc";
      when x"046a" => ROM_dataout_i <= x"78";
      when x"046b" => ROM_dataout_i <= x"cc";
      when x"046c" => ROM_dataout_i <= x"c0";
      when x"046d" => ROM_dataout_i <= x"cc";
      when x"046e" => ROM_dataout_i <= x"78";
      when x"0470" => ROM_dataout_i <= x"1c";
      when x"0471" => ROM_dataout_i <= x"0c";
      when x"0472" => ROM_dataout_i <= x"0c";
      when x"0473" => ROM_dataout_i <= x"7c";
      when x"0474" => ROM_dataout_i <= x"cc";
      when x"0475" => ROM_dataout_i <= x"cc";
      when x"0476" => ROM_dataout_i <= x"76";
      when x"047a" => ROM_dataout_i <= x"78";
      when x"047b" => ROM_dataout_i <= x"cc";
      when x"047c" => ROM_dataout_i <= x"fc";
      when x"047d" => ROM_dataout_i <= x"c0";
      when x"047e" => ROM_dataout_i <= x"78";
      when x"0480" => ROM_dataout_i <= x"38";
      when x"0481" => ROM_dataout_i <= x"6c";
      when x"0482" => ROM_dataout_i <= x"60";
      when x"0483" => ROM_dataout_i <= x"f0";
      when x"0484" => ROM_dataout_i <= x"60";
      when x"0485" => ROM_dataout_i <= x"60";
      when x"0486" => ROM_dataout_i <= x"f0";
      when x"048a" => ROM_dataout_i <= x"76";
      when x"048b" => ROM_dataout_i <= x"cc";
      when x"048c" => ROM_dataout_i <= x"cc";
      when x"048d" => ROM_dataout_i <= x"7c";
      when x"048e" => ROM_dataout_i <= x"0c";
      when x"048f" => ROM_dataout_i <= x"f8";
      when x"0490" => ROM_dataout_i <= x"e0";
      when x"0491" => ROM_dataout_i <= x"60";
      when x"0492" => ROM_dataout_i <= x"6c";
      when x"0493" => ROM_dataout_i <= x"76";
      when x"0494" => ROM_dataout_i <= x"66";
      when x"0495" => ROM_dataout_i <= x"66";
      when x"0496" => ROM_dataout_i <= x"e6";
      when x"0498" => ROM_dataout_i <= x"30";
      when x"049a" => ROM_dataout_i <= x"70";
      when x"049b" => ROM_dataout_i <= x"30";
      when x"049c" => ROM_dataout_i <= x"30";
      when x"049d" => ROM_dataout_i <= x"30";
      when x"049e" => ROM_dataout_i <= x"78";
      when x"04a0" => ROM_dataout_i <= x"0c";
      when x"04a2" => ROM_dataout_i <= x"0c";
      when x"04a3" => ROM_dataout_i <= x"0c";
      when x"04a4" => ROM_dataout_i <= x"0c";
      when x"04a5" => ROM_dataout_i <= x"cc";
      when x"04a6" => ROM_dataout_i <= x"cc";
      when x"04a7" => ROM_dataout_i <= x"78";
      when x"04a8" => ROM_dataout_i <= x"e0";
      when x"04a9" => ROM_dataout_i <= x"60";
      when x"04aa" => ROM_dataout_i <= x"66";
      when x"04ab" => ROM_dataout_i <= x"6c";
      when x"04ac" => ROM_dataout_i <= x"78";
      when x"04ad" => ROM_dataout_i <= x"6c";
      when x"04ae" => ROM_dataout_i <= x"e6";
      when x"04b0" => ROM_dataout_i <= x"70";
      when x"04b1" => ROM_dataout_i <= x"30";
      when x"04b2" => ROM_dataout_i <= x"30";
      when x"04b3" => ROM_dataout_i <= x"30";
      when x"04b4" => ROM_dataout_i <= x"30";
      when x"04b5" => ROM_dataout_i <= x"30";
      when x"04b6" => ROM_dataout_i <= x"78";
      when x"04ba" => ROM_dataout_i <= x"cc";
      when x"04bb" => ROM_dataout_i <= x"fe";
      when x"04bc" => ROM_dataout_i <= x"fe";
      when x"04bd" => ROM_dataout_i <= x"d6";
      when x"04be" => ROM_dataout_i <= x"c6";
      when x"04c2" => ROM_dataout_i <= x"f8";
      when x"04c3" => ROM_dataout_i <= x"cc";
      when x"04c4" => ROM_dataout_i <= x"cc";
      when x"04c5" => ROM_dataout_i <= x"cc";
      when x"04c6" => ROM_dataout_i <= x"cc";
      when x"04ca" => ROM_dataout_i <= x"78";
      when x"04cb" => ROM_dataout_i <= x"cc";
      when x"04cc" => ROM_dataout_i <= x"cc";
      when x"04cd" => ROM_dataout_i <= x"cc";
      when x"04ce" => ROM_dataout_i <= x"78";
      when x"04d2" => ROM_dataout_i <= x"dc";
      when x"04d3" => ROM_dataout_i <= x"66";
      when x"04d4" => ROM_dataout_i <= x"66";
      when x"04d5" => ROM_dataout_i <= x"7c";
      when x"04d6" => ROM_dataout_i <= x"60";
      when x"04d7" => ROM_dataout_i <= x"f0";
      when x"04da" => ROM_dataout_i <= x"76";
      when x"04db" => ROM_dataout_i <= x"cc";
      when x"04dc" => ROM_dataout_i <= x"cc";
      when x"04dd" => ROM_dataout_i <= x"7c";
      when x"04de" => ROM_dataout_i <= x"0c";
      when x"04df" => ROM_dataout_i <= x"1e";
      when x"04e2" => ROM_dataout_i <= x"dc";
      when x"04e3" => ROM_dataout_i <= x"76";
      when x"04e4" => ROM_dataout_i <= x"66";
      when x"04e5" => ROM_dataout_i <= x"60";
      when x"04e6" => ROM_dataout_i <= x"f0";
      when x"04ea" => ROM_dataout_i <= x"7c";
      when x"04eb" => ROM_dataout_i <= x"c0";
      when x"04ec" => ROM_dataout_i <= x"78";
      when x"04ed" => ROM_dataout_i <= x"0c";
      when x"04ee" => ROM_dataout_i <= x"f8";
      when x"04f0" => ROM_dataout_i <= x"10";
      when x"04f1" => ROM_dataout_i <= x"30";
      when x"04f2" => ROM_dataout_i <= x"7c";
      when x"04f3" => ROM_dataout_i <= x"30";
      when x"04f4" => ROM_dataout_i <= x"30";
      when x"04f5" => ROM_dataout_i <= x"34";
      when x"04f6" => ROM_dataout_i <= x"18";
      when x"04fa" => ROM_dataout_i <= x"cc";
      when x"04fb" => ROM_dataout_i <= x"cc";
      when x"04fc" => ROM_dataout_i <= x"cc";
      when x"04fd" => ROM_dataout_i <= x"cc";
      when x"04fe" => ROM_dataout_i <= x"76";
      when x"0502" => ROM_dataout_i <= x"cc";
      when x"0503" => ROM_dataout_i <= x"cc";
      when x"0504" => ROM_dataout_i <= x"cc";
      when x"0505" => ROM_dataout_i <= x"78";
      when x"0506" => ROM_dataout_i <= x"30";
      when x"050a" => ROM_dataout_i <= x"c6";
      when x"050b" => ROM_dataout_i <= x"d6";
      when x"050c" => ROM_dataout_i <= x"fe";
      when x"050d" => ROM_dataout_i <= x"fe";
      when x"050e" => ROM_dataout_i <= x"6c";
      when x"0512" => ROM_dataout_i <= x"c6";
      when x"0513" => ROM_dataout_i <= x"6c";
      when x"0514" => ROM_dataout_i <= x"38";
      when x"0515" => ROM_dataout_i <= x"6c";
      when x"0516" => ROM_dataout_i <= x"c6";
      when x"051a" => ROM_dataout_i <= x"cc";
      when x"051b" => ROM_dataout_i <= x"cc";
      when x"051c" => ROM_dataout_i <= x"cc";
      when x"051d" => ROM_dataout_i <= x"7c";
      when x"051e" => ROM_dataout_i <= x"0c";
      when x"051f" => ROM_dataout_i <= x"f8";
      when x"0522" => ROM_dataout_i <= x"fc";
      when x"0523" => ROM_dataout_i <= x"98";
      when x"0524" => ROM_dataout_i <= x"30";
      when x"0525" => ROM_dataout_i <= x"64";
      when x"0526" => ROM_dataout_i <= x"fc";
      when x"0528" => ROM_dataout_i <= x"1c";
      when x"0529" => ROM_dataout_i <= x"30";
      when x"052a" => ROM_dataout_i <= x"30";
      when x"052b" => ROM_dataout_i <= x"e0";
      when x"052c" => ROM_dataout_i <= x"30";
      when x"052d" => ROM_dataout_i <= x"30";
      when x"052e" => ROM_dataout_i <= x"1c";
      when x"0530" => ROM_dataout_i <= x"18";
      when x"0531" => ROM_dataout_i <= x"18";
      when x"0532" => ROM_dataout_i <= x"18";
      when x"0534" => ROM_dataout_i <= x"18";
      when x"0535" => ROM_dataout_i <= x"18";
      when x"0536" => ROM_dataout_i <= x"18";
      when x"0538" => ROM_dataout_i <= x"e0";
      when x"0539" => ROM_dataout_i <= x"30";
      when x"053a" => ROM_dataout_i <= x"30";
      when x"053b" => ROM_dataout_i <= x"1c";
      when x"053c" => ROM_dataout_i <= x"30";
      when x"053d" => ROM_dataout_i <= x"30";
      when x"053e" => ROM_dataout_i <= x"e0";
      when x"0540" => ROM_dataout_i <= x"76";
      when x"0541" => ROM_dataout_i <= x"dc";
      when x"0549" => ROM_dataout_i <= x"10";
      when x"054a" => ROM_dataout_i <= x"38";
      when x"054b" => ROM_dataout_i <= x"6c";
      when x"054c" => ROM_dataout_i <= x"c6";
      when x"054d" => ROM_dataout_i <= x"fe";
      when x"0550" => ROM_dataout_i <= x"3c";
      when x"0551" => ROM_dataout_i <= x"66";
      when x"0552" => ROM_dataout_i <= x"c0";
      when x"0553" => ROM_dataout_i <= x"c0";
      when x"0554" => ROM_dataout_i <= x"66";
      when x"0555" => ROM_dataout_i <= x"3c";
      when x"0556" => ROM_dataout_i <= x"08";
      when x"0557" => ROM_dataout_i <= x"18";
      when x"0558" => ROM_dataout_i <= x"28";
      when x"055a" => ROM_dataout_i <= x"cc";
      when x"055b" => ROM_dataout_i <= x"cc";
      when x"055c" => ROM_dataout_i <= x"cc";
      when x"055d" => ROM_dataout_i <= x"cc";
      when x"055e" => ROM_dataout_i <= x"76";
      when x"0560" => ROM_dataout_i <= x"08";
      when x"0561" => ROM_dataout_i <= x"10";
      when x"0562" => ROM_dataout_i <= x"78";
      when x"0563" => ROM_dataout_i <= x"cc";
      when x"0564" => ROM_dataout_i <= x"fc";
      when x"0565" => ROM_dataout_i <= x"c0";
      when x"0566" => ROM_dataout_i <= x"78";
      when x"0568" => ROM_dataout_i <= x"10";
      when x"0569" => ROM_dataout_i <= x"28";
      when x"056a" => ROM_dataout_i <= x"78";
      when x"056b" => ROM_dataout_i <= x"0c";
      when x"056c" => ROM_dataout_i <= x"7c";
      when x"056d" => ROM_dataout_i <= x"cc";
      when x"056e" => ROM_dataout_i <= x"76";
      when x"0570" => ROM_dataout_i <= x"28";
      when x"0572" => ROM_dataout_i <= x"78";
      when x"0573" => ROM_dataout_i <= x"0c";
      when x"0574" => ROM_dataout_i <= x"7c";
      when x"0575" => ROM_dataout_i <= x"cc";
      when x"0576" => ROM_dataout_i <= x"76";
      when x"0578" => ROM_dataout_i <= x"20";
      when x"0579" => ROM_dataout_i <= x"10";
      when x"057a" => ROM_dataout_i <= x"78";
      when x"057b" => ROM_dataout_i <= x"0c";
      when x"057c" => ROM_dataout_i <= x"7c";
      when x"057d" => ROM_dataout_i <= x"cc";
      when x"057e" => ROM_dataout_i <= x"76";
      when x"0580" => ROM_dataout_i <= x"18";
      when x"0581" => ROM_dataout_i <= x"18";
      when x"0582" => ROM_dataout_i <= x"78";
      when x"0583" => ROM_dataout_i <= x"0c";
      when x"0584" => ROM_dataout_i <= x"7c";
      when x"0585" => ROM_dataout_i <= x"cc";
      when x"0586" => ROM_dataout_i <= x"76";
      when x"0589" => ROM_dataout_i <= x"78";
      when x"058a" => ROM_dataout_i <= x"cc";
      when x"058b" => ROM_dataout_i <= x"c0";
      when x"058c" => ROM_dataout_i <= x"cc";
      when x"058d" => ROM_dataout_i <= x"78";
      when x"058e" => ROM_dataout_i <= x"10";
      when x"058f" => ROM_dataout_i <= x"30";
      when x"0590" => ROM_dataout_i <= x"10";
      when x"0591" => ROM_dataout_i <= x"28";
      when x"0592" => ROM_dataout_i <= x"78";
      when x"0593" => ROM_dataout_i <= x"cc";
      when x"0594" => ROM_dataout_i <= x"fc";
      when x"0595" => ROM_dataout_i <= x"c0";
      when x"0596" => ROM_dataout_i <= x"78";
      when x"0598" => ROM_dataout_i <= x"28";
      when x"059a" => ROM_dataout_i <= x"78";
      when x"059b" => ROM_dataout_i <= x"cc";
      when x"059c" => ROM_dataout_i <= x"fc";
      when x"059d" => ROM_dataout_i <= x"c0";
      when x"059e" => ROM_dataout_i <= x"78";
      when x"05a0" => ROM_dataout_i <= x"20";
      when x"05a1" => ROM_dataout_i <= x"10";
      when x"05a2" => ROM_dataout_i <= x"78";
      when x"05a3" => ROM_dataout_i <= x"cc";
      when x"05a4" => ROM_dataout_i <= x"fc";
      when x"05a5" => ROM_dataout_i <= x"c0";
      when x"05a6" => ROM_dataout_i <= x"78";
      when x"05a8" => ROM_dataout_i <= x"28";
      when x"05aa" => ROM_dataout_i <= x"70";
      when x"05ab" => ROM_dataout_i <= x"30";
      when x"05ac" => ROM_dataout_i <= x"30";
      when x"05ad" => ROM_dataout_i <= x"30";
      when x"05ae" => ROM_dataout_i <= x"78";
      when x"05b0" => ROM_dataout_i <= x"10";
      when x"05b1" => ROM_dataout_i <= x"28";
      when x"05b2" => ROM_dataout_i <= x"70";
      when x"05b3" => ROM_dataout_i <= x"30";
      when x"05b4" => ROM_dataout_i <= x"30";
      when x"05b5" => ROM_dataout_i <= x"30";
      when x"05b6" => ROM_dataout_i <= x"78";
      when x"05b8" => ROM_dataout_i <= x"10";
      when x"05b9" => ROM_dataout_i <= x"08";
      when x"05ba" => ROM_dataout_i <= x"70";
      when x"05bb" => ROM_dataout_i <= x"30";
      when x"05bc" => ROM_dataout_i <= x"30";
      when x"05bd" => ROM_dataout_i <= x"30";
      when x"05be" => ROM_dataout_i <= x"78";
      when x"05c0" => ROM_dataout_i <= x"28";
      when x"05c1" => ROM_dataout_i <= x"30";
      when x"05c2" => ROM_dataout_i <= x"78";
      when x"05c3" => ROM_dataout_i <= x"cc";
      when x"05c4" => ROM_dataout_i <= x"fc";
      when x"05c5" => ROM_dataout_i <= x"cc";
      when x"05c6" => ROM_dataout_i <= x"cc";
      when x"05c8" => ROM_dataout_i <= x"30";
      when x"05c9" => ROM_dataout_i <= x"48";
      when x"05ca" => ROM_dataout_i <= x"30";
      when x"05cb" => ROM_dataout_i <= x"cc";
      when x"05cc" => ROM_dataout_i <= x"fc";
      when x"05cd" => ROM_dataout_i <= x"cc";
      when x"05ce" => ROM_dataout_i <= x"cc";
      when x"05d0" => ROM_dataout_i <= x"08";
      when x"05d1" => ROM_dataout_i <= x"10";
      when x"05d2" => ROM_dataout_i <= x"7e";
      when x"05d3" => ROM_dataout_i <= x"60";
      when x"05d4" => ROM_dataout_i <= x"78";
      when x"05d5" => ROM_dataout_i <= x"60";
      when x"05d6" => ROM_dataout_i <= x"7e";
      when x"05da" => ROM_dataout_i <= x"6c";
      when x"05db" => ROM_dataout_i <= x"12";
      when x"05dc" => ROM_dataout_i <= x"7e";
      when x"05dd" => ROM_dataout_i <= x"90";
      when x"05de" => ROM_dataout_i <= x"7e";
      when x"05e0" => ROM_dataout_i <= x"3e";
      when x"05e1" => ROM_dataout_i <= x"50";
      when x"05e2" => ROM_dataout_i <= x"90";
      when x"05e3" => ROM_dataout_i <= x"9c";
      when x"05e4" => ROM_dataout_i <= x"f0";
      when x"05e5" => ROM_dataout_i <= x"90";
      when x"05e6" => ROM_dataout_i <= x"9e";
      when x"05e8" => ROM_dataout_i <= x"10";
      when x"05e9" => ROM_dataout_i <= x"28";
      when x"05ea" => ROM_dataout_i <= x"78";
      when x"05eb" => ROM_dataout_i <= x"cc";
      when x"05ec" => ROM_dataout_i <= x"cc";
      when x"05ed" => ROM_dataout_i <= x"cc";
      when x"05ee" => ROM_dataout_i <= x"78";
      when x"05f0" => ROM_dataout_i <= x"28";
      when x"05f2" => ROM_dataout_i <= x"78";
      when x"05f3" => ROM_dataout_i <= x"cc";
      when x"05f4" => ROM_dataout_i <= x"cc";
      when x"05f5" => ROM_dataout_i <= x"cc";
      when x"05f6" => ROM_dataout_i <= x"78";
      when x"05f8" => ROM_dataout_i <= x"20";
      when x"05f9" => ROM_dataout_i <= x"10";
      when x"05fa" => ROM_dataout_i <= x"78";
      when x"05fb" => ROM_dataout_i <= x"cc";
      when x"05fc" => ROM_dataout_i <= x"cc";
      when x"05fd" => ROM_dataout_i <= x"cc";
      when x"05fe" => ROM_dataout_i <= x"78";
      when x"0600" => ROM_dataout_i <= x"10";
      when x"0601" => ROM_dataout_i <= x"28";
      when x"0602" => ROM_dataout_i <= x"cc";
      when x"0603" => ROM_dataout_i <= x"cc";
      when x"0604" => ROM_dataout_i <= x"cc";
      when x"0605" => ROM_dataout_i <= x"cc";
      when x"0606" => ROM_dataout_i <= x"76";
      when x"0608" => ROM_dataout_i <= x"20";
      when x"0609" => ROM_dataout_i <= x"10";
      when x"060a" => ROM_dataout_i <= x"cc";
      when x"060b" => ROM_dataout_i <= x"cc";
      when x"060c" => ROM_dataout_i <= x"cc";
      when x"060d" => ROM_dataout_i <= x"cc";
      when x"060e" => ROM_dataout_i <= x"76";
      when x"0610" => ROM_dataout_i <= x"28";
      when x"0612" => ROM_dataout_i <= x"cc";
      when x"0613" => ROM_dataout_i <= x"cc";
      when x"0614" => ROM_dataout_i <= x"cc";
      when x"0615" => ROM_dataout_i <= x"7c";
      when x"0616" => ROM_dataout_i <= x"0c";
      when x"0617" => ROM_dataout_i <= x"f8";
      when x"0618" => ROM_dataout_i <= x"28";
      when x"0619" => ROM_dataout_i <= x"7c";
      when x"061a" => ROM_dataout_i <= x"c6";
      when x"061b" => ROM_dataout_i <= x"c6";
      when x"061c" => ROM_dataout_i <= x"c6";
      when x"061d" => ROM_dataout_i <= x"c6";
      when x"061e" => ROM_dataout_i <= x"7c";
      when x"0620" => ROM_dataout_i <= x"28";
      when x"0621" => ROM_dataout_i <= x"c6";
      when x"0622" => ROM_dataout_i <= x"c6";
      when x"0623" => ROM_dataout_i <= x"c6";
      when x"0624" => ROM_dataout_i <= x"c6";
      when x"0625" => ROM_dataout_i <= x"c6";
      when x"0626" => ROM_dataout_i <= x"7c";
      when x"0629" => ROM_dataout_i <= x"10";
      when x"062a" => ROM_dataout_i <= x"78";
      when x"062b" => ROM_dataout_i <= x"cc";
      when x"062c" => ROM_dataout_i <= x"c0";
      when x"062d" => ROM_dataout_i <= x"cc";
      when x"062e" => ROM_dataout_i <= x"78";
      when x"062f" => ROM_dataout_i <= x"10";
      when x"0630" => ROM_dataout_i <= x"38";
      when x"0631" => ROM_dataout_i <= x"44";
      when x"0632" => ROM_dataout_i <= x"40";
      when x"0633" => ROM_dataout_i <= x"f0";
      when x"0634" => ROM_dataout_i <= x"40";
      when x"0635" => ROM_dataout_i <= x"40";
      when x"0636" => ROM_dataout_i <= x"fe";
      when x"0638" => ROM_dataout_i <= x"c3";
      when x"0639" => ROM_dataout_i <= x"66";
      when x"063a" => ROM_dataout_i <= x"3c";
      when x"063b" => ROM_dataout_i <= x"7e";
      when x"063c" => ROM_dataout_i <= x"18";
      when x"063d" => ROM_dataout_i <= x"7e";
      when x"063e" => ROM_dataout_i <= x"18";
      when x"0640" => ROM_dataout_i <= x"fc";
      when x"0641" => ROM_dataout_i <= x"66";
      when x"0642" => ROM_dataout_i <= x"66";
      when x"0643" => ROM_dataout_i <= x"7c";
      when x"0644" => ROM_dataout_i <= x"60";
      when x"0645" => ROM_dataout_i <= x"60";
      when x"0646" => ROM_dataout_i <= x"f0";
      when x"0648" => ROM_dataout_i <= x"1c";
      when x"0649" => ROM_dataout_i <= x"30";
      when x"064a" => ROM_dataout_i <= x"fc";
      when x"064b" => ROM_dataout_i <= x"30";
      when x"064c" => ROM_dataout_i <= x"30";
      when x"064d" => ROM_dataout_i <= x"30";
      when x"064e" => ROM_dataout_i <= x"30";
      when x"064f" => ROM_dataout_i <= x"e0";
      when x"0650" => ROM_dataout_i <= x"08";
      when x"0651" => ROM_dataout_i <= x"10";
      when x"0652" => ROM_dataout_i <= x"78";
      when x"0653" => ROM_dataout_i <= x"0c";
      when x"0654" => ROM_dataout_i <= x"7c";
      when x"0655" => ROM_dataout_i <= x"cc";
      when x"0656" => ROM_dataout_i <= x"76";
      when x"0658" => ROM_dataout_i <= x"10";
      when x"0659" => ROM_dataout_i <= x"20";
      when x"065a" => ROM_dataout_i <= x"70";
      when x"065b" => ROM_dataout_i <= x"30";
      when x"065c" => ROM_dataout_i <= x"30";
      when x"065d" => ROM_dataout_i <= x"30";
      when x"065e" => ROM_dataout_i <= x"78";
      when x"0660" => ROM_dataout_i <= x"10";
      when x"0661" => ROM_dataout_i <= x"20";
      when x"0662" => ROM_dataout_i <= x"78";
      when x"0663" => ROM_dataout_i <= x"cc";
      when x"0664" => ROM_dataout_i <= x"cc";
      when x"0665" => ROM_dataout_i <= x"cc";
      when x"0666" => ROM_dataout_i <= x"78";
      when x"0668" => ROM_dataout_i <= x"10";
      when x"0669" => ROM_dataout_i <= x"20";
      when x"066a" => ROM_dataout_i <= x"cc";
      when x"066b" => ROM_dataout_i <= x"cc";
      when x"066c" => ROM_dataout_i <= x"cc";
      when x"066d" => ROM_dataout_i <= x"cc";
      when x"066e" => ROM_dataout_i <= x"76";
      when x"0670" => ROM_dataout_i <= x"32";
      when x"0671" => ROM_dataout_i <= x"4c";
      when x"0672" => ROM_dataout_i <= x"f8";
      when x"0673" => ROM_dataout_i <= x"cc";
      when x"0674" => ROM_dataout_i <= x"cc";
      when x"0675" => ROM_dataout_i <= x"cc";
      when x"0676" => ROM_dataout_i <= x"cc";
      when x"0678" => ROM_dataout_i <= x"32";
      when x"0679" => ROM_dataout_i <= x"4c";
      when x"067a" => ROM_dataout_i <= x"c6";
      when x"067b" => ROM_dataout_i <= x"e6";
      when x"067c" => ROM_dataout_i <= x"d6";
      when x"067d" => ROM_dataout_i <= x"ce";
      when x"067e" => ROM_dataout_i <= x"c6";
      when x"0681" => ROM_dataout_i <= x"38";
      when x"0682" => ROM_dataout_i <= x"0c";
      when x"0683" => ROM_dataout_i <= x"3c";
      when x"0684" => ROM_dataout_i <= x"6c";
      when x"0685" => ROM_dataout_i <= x"36";
      when x"0689" => ROM_dataout_i <= x"38";
      when x"068a" => ROM_dataout_i <= x"44";
      when x"068b" => ROM_dataout_i <= x"44";
      when x"068c" => ROM_dataout_i <= x"38";
      when x"0690" => ROM_dataout_i <= x"18";
      when x"0692" => ROM_dataout_i <= x"18";
      when x"0693" => ROM_dataout_i <= x"30";
      when x"0694" => ROM_dataout_i <= x"60";
      when x"0695" => ROM_dataout_i <= x"66";
      when x"0696" => ROM_dataout_i <= x"3c";
      when x"069a" => ROM_dataout_i <= x"fe";
      when x"069b" => ROM_dataout_i <= x"80";
      when x"069c" => ROM_dataout_i <= x"80";
      when x"06a2" => ROM_dataout_i <= x"fe";
      when x"06a3" => ROM_dataout_i <= x"02";
      when x"06a4" => ROM_dataout_i <= x"02";
      when x"06a8" => ROM_dataout_i <= x"42";
      when x"06a9" => ROM_dataout_i <= x"44";
      when x"06aa" => ROM_dataout_i <= x"48";
      when x"06ab" => ROM_dataout_i <= x"56";
      when x"06ac" => ROM_dataout_i <= x"29";
      when x"06ad" => ROM_dataout_i <= x"46";
      when x"06ae" => ROM_dataout_i <= x"88";
      when x"06af" => ROM_dataout_i <= x"1f";
      when x"06b0" => ROM_dataout_i <= x"42";
      when x"06b1" => ROM_dataout_i <= x"44";
      when x"06b2" => ROM_dataout_i <= x"48";
      when x"06b3" => ROM_dataout_i <= x"56";
      when x"06b4" => ROM_dataout_i <= x"2a";
      when x"06b5" => ROM_dataout_i <= x"5f";
      when x"06b6" => ROM_dataout_i <= x"82";
      when x"06b7" => ROM_dataout_i <= x"07";
      when x"06b8" => ROM_dataout_i <= x"30";
      when x"06ba" => ROM_dataout_i <= x"30";
      when x"06bb" => ROM_dataout_i <= x"30";
      when x"06bc" => ROM_dataout_i <= x"30";
      when x"06bd" => ROM_dataout_i <= x"30";
      when x"06be" => ROM_dataout_i <= x"30";
      when x"06c1" => ROM_dataout_i <= x"24";
      when x"06c2" => ROM_dataout_i <= x"48";
      when x"06c3" => ROM_dataout_i <= x"90";
      when x"06c4" => ROM_dataout_i <= x"48";
      when x"06c5" => ROM_dataout_i <= x"24";
      when x"06c9" => ROM_dataout_i <= x"48";
      when x"06ca" => ROM_dataout_i <= x"24";
      when x"06cb" => ROM_dataout_i <= x"12";
      when x"06cc" => ROM_dataout_i <= x"24";
      when x"06cd" => ROM_dataout_i <= x"48";
      when x"06d0" => ROM_dataout_i <= x"88";
      when x"06d1" => ROM_dataout_i <= x"22";
      when x"06d2" => ROM_dataout_i <= x"88";
      when x"06d3" => ROM_dataout_i <= x"22";
      when x"06d4" => ROM_dataout_i <= x"88";
      when x"06d6" => ROM_dataout_i <= x"88";
      when x"06d7" => ROM_dataout_i <= x"22";
      when x"06d8" => ROM_dataout_i <= x"aa";
      when x"06d9" => ROM_dataout_i <= x"55";
      when x"06da" => ROM_dataout_i <= x"aa";
      when x"06db" => ROM_dataout_i <= x"55";
      when x"06dc" => ROM_dataout_i <= x"aa";
      when x"06de" => ROM_dataout_i <= x"aa";
      when x"06df" => ROM_dataout_i <= x"55";
      when x"06e0" => ROM_dataout_i <= x"77";
      when x"06e1" => ROM_dataout_i <= x"dd";
      when x"06e2" => ROM_dataout_i <= x"77";
      when x"06e3" => ROM_dataout_i <= x"dd";
      when x"06e4" => ROM_dataout_i <= x"77";
      when x"06e5" => ROM_dataout_i <= x"ff";
      when x"06e6" => ROM_dataout_i <= x"77";
      when x"06e7" => ROM_dataout_i <= x"dd";
      when x"06e8" => ROM_dataout_i <= x"10";
      when x"06e9" => ROM_dataout_i <= x"10";
      when x"06ea" => ROM_dataout_i <= x"10";
      when x"06eb" => ROM_dataout_i <= x"10";
      when x"06ec" => ROM_dataout_i <= x"10";
      when x"06ed" => ROM_dataout_i <= x"10";
      when x"06ee" => ROM_dataout_i <= x"10";
      when x"06ef" => ROM_dataout_i <= x"10";
      when x"06f0" => ROM_dataout_i <= x"10";
      when x"06f1" => ROM_dataout_i <= x"10";
      when x"06f2" => ROM_dataout_i <= x"10";
      when x"06f3" => ROM_dataout_i <= x"f0";
      when x"06f4" => ROM_dataout_i <= x"10";
      when x"06f5" => ROM_dataout_i <= x"10";
      when x"06f6" => ROM_dataout_i <= x"10";
      when x"06f7" => ROM_dataout_i <= x"10";
      when x"06f8" => ROM_dataout_i <= x"10";
      when x"06f9" => ROM_dataout_i <= x"10";
      when x"06fa" => ROM_dataout_i <= x"f0";
      when x"06fb" => ROM_dataout_i <= x"10";
      when x"06fc" => ROM_dataout_i <= x"f0";
      when x"06fd" => ROM_dataout_i <= x"10";
      when x"06fe" => ROM_dataout_i <= x"10";
      when x"06ff" => ROM_dataout_i <= x"10";
      when x"0700" => ROM_dataout_i <= x"28";
      when x"0701" => ROM_dataout_i <= x"28";
      when x"0702" => ROM_dataout_i <= x"28";
      when x"0703" => ROM_dataout_i <= x"e8";
      when x"0704" => ROM_dataout_i <= x"28";
      when x"0705" => ROM_dataout_i <= x"28";
      when x"0706" => ROM_dataout_i <= x"28";
      when x"0707" => ROM_dataout_i <= x"28";
      when x"070b" => ROM_dataout_i <= x"f8";
      when x"070c" => ROM_dataout_i <= x"28";
      when x"070d" => ROM_dataout_i <= x"28";
      when x"070e" => ROM_dataout_i <= x"28";
      when x"070f" => ROM_dataout_i <= x"28";
      when x"0712" => ROM_dataout_i <= x"f0";
      when x"0713" => ROM_dataout_i <= x"10";
      when x"0714" => ROM_dataout_i <= x"f0";
      when x"0715" => ROM_dataout_i <= x"10";
      when x"0716" => ROM_dataout_i <= x"10";
      when x"0717" => ROM_dataout_i <= x"10";
      when x"0718" => ROM_dataout_i <= x"28";
      when x"0719" => ROM_dataout_i <= x"28";
      when x"071a" => ROM_dataout_i <= x"e8";
      when x"071b" => ROM_dataout_i <= x"08";
      when x"071c" => ROM_dataout_i <= x"e8";
      when x"071d" => ROM_dataout_i <= x"28";
      when x"071e" => ROM_dataout_i <= x"28";
      when x"071f" => ROM_dataout_i <= x"28";
      when x"0720" => ROM_dataout_i <= x"28";
      when x"0721" => ROM_dataout_i <= x"28";
      when x"0722" => ROM_dataout_i <= x"28";
      when x"0723" => ROM_dataout_i <= x"28";
      when x"0724" => ROM_dataout_i <= x"28";
      when x"0725" => ROM_dataout_i <= x"28";
      when x"0726" => ROM_dataout_i <= x"28";
      when x"0727" => ROM_dataout_i <= x"28";
      when x"072a" => ROM_dataout_i <= x"f8";
      when x"072b" => ROM_dataout_i <= x"08";
      when x"072c" => ROM_dataout_i <= x"e8";
      when x"072d" => ROM_dataout_i <= x"28";
      when x"072e" => ROM_dataout_i <= x"28";
      when x"072f" => ROM_dataout_i <= x"28";
      when x"0730" => ROM_dataout_i <= x"28";
      when x"0731" => ROM_dataout_i <= x"28";
      when x"0732" => ROM_dataout_i <= x"e8";
      when x"0733" => ROM_dataout_i <= x"08";
      when x"0734" => ROM_dataout_i <= x"f8";
      when x"0738" => ROM_dataout_i <= x"28";
      when x"0739" => ROM_dataout_i <= x"28";
      when x"073a" => ROM_dataout_i <= x"28";
      when x"073b" => ROM_dataout_i <= x"f8";
      when x"0740" => ROM_dataout_i <= x"10";
      when x"0741" => ROM_dataout_i <= x"10";
      when x"0742" => ROM_dataout_i <= x"f0";
      when x"0743" => ROM_dataout_i <= x"10";
      when x"0744" => ROM_dataout_i <= x"f0";
      when x"074b" => ROM_dataout_i <= x"f0";
      when x"074c" => ROM_dataout_i <= x"10";
      when x"074d" => ROM_dataout_i <= x"10";
      when x"074e" => ROM_dataout_i <= x"10";
      when x"074f" => ROM_dataout_i <= x"10";
      when x"0750" => ROM_dataout_i <= x"10";
      when x"0751" => ROM_dataout_i <= x"10";
      when x"0752" => ROM_dataout_i <= x"10";
      when x"0753" => ROM_dataout_i <= x"1f";
      when x"0758" => ROM_dataout_i <= x"10";
      when x"0759" => ROM_dataout_i <= x"10";
      when x"075a" => ROM_dataout_i <= x"10";
      when x"075b" => ROM_dataout_i <= x"ff";
      when x"0763" => ROM_dataout_i <= x"ff";
      when x"0764" => ROM_dataout_i <= x"10";
      when x"0765" => ROM_dataout_i <= x"10";
      when x"0766" => ROM_dataout_i <= x"10";
      when x"0767" => ROM_dataout_i <= x"10";
      when x"0768" => ROM_dataout_i <= x"10";
      when x"0769" => ROM_dataout_i <= x"10";
      when x"076a" => ROM_dataout_i <= x"10";
      when x"076b" => ROM_dataout_i <= x"1f";
      when x"076c" => ROM_dataout_i <= x"10";
      when x"076d" => ROM_dataout_i <= x"10";
      when x"076e" => ROM_dataout_i <= x"10";
      when x"076f" => ROM_dataout_i <= x"10";
      when x"0773" => ROM_dataout_i <= x"ff";
      when x"0778" => ROM_dataout_i <= x"10";
      when x"0779" => ROM_dataout_i <= x"10";
      when x"077a" => ROM_dataout_i <= x"10";
      when x"077b" => ROM_dataout_i <= x"ff";
      when x"077c" => ROM_dataout_i <= x"10";
      when x"077d" => ROM_dataout_i <= x"10";
      when x"077e" => ROM_dataout_i <= x"10";
      when x"077f" => ROM_dataout_i <= x"10";
      when x"0780" => ROM_dataout_i <= x"10";
      when x"0781" => ROM_dataout_i <= x"10";
      when x"0782" => ROM_dataout_i <= x"1f";
      when x"0783" => ROM_dataout_i <= x"10";
      when x"0784" => ROM_dataout_i <= x"1f";
      when x"0785" => ROM_dataout_i <= x"10";
      when x"0786" => ROM_dataout_i <= x"10";
      when x"0787" => ROM_dataout_i <= x"10";
      when x"0788" => ROM_dataout_i <= x"28";
      when x"0789" => ROM_dataout_i <= x"28";
      when x"078a" => ROM_dataout_i <= x"28";
      when x"078b" => ROM_dataout_i <= x"2f";
      when x"078c" => ROM_dataout_i <= x"28";
      when x"078d" => ROM_dataout_i <= x"28";
      when x"078e" => ROM_dataout_i <= x"28";
      when x"078f" => ROM_dataout_i <= x"28";
      when x"0790" => ROM_dataout_i <= x"28";
      when x"0791" => ROM_dataout_i <= x"28";
      when x"0792" => ROM_dataout_i <= x"2f";
      when x"0793" => ROM_dataout_i <= x"20";
      when x"0794" => ROM_dataout_i <= x"3f";
      when x"079a" => ROM_dataout_i <= x"3f";
      when x"079b" => ROM_dataout_i <= x"20";
      when x"079c" => ROM_dataout_i <= x"2f";
      when x"079d" => ROM_dataout_i <= x"28";
      when x"079e" => ROM_dataout_i <= x"28";
      when x"079f" => ROM_dataout_i <= x"28";
      when x"07a0" => ROM_dataout_i <= x"28";
      when x"07a1" => ROM_dataout_i <= x"28";
      when x"07a2" => ROM_dataout_i <= x"ef";
      when x"07a4" => ROM_dataout_i <= x"ff";
      when x"07aa" => ROM_dataout_i <= x"ff";
      when x"07ac" => ROM_dataout_i <= x"ef";
      when x"07ad" => ROM_dataout_i <= x"28";
      when x"07ae" => ROM_dataout_i <= x"28";
      when x"07af" => ROM_dataout_i <= x"28";
      when x"07b0" => ROM_dataout_i <= x"28";
      when x"07b1" => ROM_dataout_i <= x"28";
      when x"07b2" => ROM_dataout_i <= x"2f";
      when x"07b3" => ROM_dataout_i <= x"20";
      when x"07b4" => ROM_dataout_i <= x"2f";
      when x"07b5" => ROM_dataout_i <= x"28";
      when x"07b6" => ROM_dataout_i <= x"28";
      when x"07b7" => ROM_dataout_i <= x"28";
      when x"07ba" => ROM_dataout_i <= x"ff";
      when x"07bc" => ROM_dataout_i <= x"ff";
      when x"07c0" => ROM_dataout_i <= x"28";
      when x"07c1" => ROM_dataout_i <= x"28";
      when x"07c2" => ROM_dataout_i <= x"ef";
      when x"07c4" => ROM_dataout_i <= x"ef";
      when x"07c5" => ROM_dataout_i <= x"28";
      when x"07c6" => ROM_dataout_i <= x"28";
      when x"07c7" => ROM_dataout_i <= x"28";
      when x"07c8" => ROM_dataout_i <= x"10";
      when x"07c9" => ROM_dataout_i <= x"10";
      when x"07ca" => ROM_dataout_i <= x"ff";
      when x"07cc" => ROM_dataout_i <= x"ff";
      when x"07d0" => ROM_dataout_i <= x"28";
      when x"07d1" => ROM_dataout_i <= x"28";
      when x"07d2" => ROM_dataout_i <= x"28";
      when x"07d3" => ROM_dataout_i <= x"ff";
      when x"07da" => ROM_dataout_i <= x"ff";
      when x"07dc" => ROM_dataout_i <= x"ff";
      when x"07dd" => ROM_dataout_i <= x"10";
      when x"07de" => ROM_dataout_i <= x"10";
      when x"07df" => ROM_dataout_i <= x"10";
      when x"07e3" => ROM_dataout_i <= x"ff";
      when x"07e4" => ROM_dataout_i <= x"28";
      when x"07e5" => ROM_dataout_i <= x"28";
      when x"07e6" => ROM_dataout_i <= x"28";
      when x"07e7" => ROM_dataout_i <= x"28";
      when x"07e8" => ROM_dataout_i <= x"28";
      when x"07e9" => ROM_dataout_i <= x"28";
      when x"07ea" => ROM_dataout_i <= x"28";
      when x"07eb" => ROM_dataout_i <= x"3f";
      when x"07f0" => ROM_dataout_i <= x"10";
      when x"07f1" => ROM_dataout_i <= x"10";
      when x"07f2" => ROM_dataout_i <= x"1f";
      when x"07f3" => ROM_dataout_i <= x"10";
      when x"07f4" => ROM_dataout_i <= x"1f";
      when x"07fa" => ROM_dataout_i <= x"1f";
      when x"07fb" => ROM_dataout_i <= x"10";
      when x"07fc" => ROM_dataout_i <= x"1f";
      when x"07fd" => ROM_dataout_i <= x"10";
      when x"07fe" => ROM_dataout_i <= x"10";
      when x"07ff" => ROM_dataout_i <= x"10";
      when x"0803" => ROM_dataout_i <= x"3f";
      when x"0804" => ROM_dataout_i <= x"28";
      when x"0805" => ROM_dataout_i <= x"28";
      when x"0806" => ROM_dataout_i <= x"28";
      when x"0807" => ROM_dataout_i <= x"28";
      when x"0808" => ROM_dataout_i <= x"28";
      when x"0809" => ROM_dataout_i <= x"28";
      when x"080a" => ROM_dataout_i <= x"28";
      when x"080b" => ROM_dataout_i <= x"ff";
      when x"080c" => ROM_dataout_i <= x"28";
      when x"080d" => ROM_dataout_i <= x"28";
      when x"080e" => ROM_dataout_i <= x"28";
      when x"080f" => ROM_dataout_i <= x"28";
      when x"0810" => ROM_dataout_i <= x"10";
      when x"0811" => ROM_dataout_i <= x"10";
      when x"0812" => ROM_dataout_i <= x"ff";
      when x"0813" => ROM_dataout_i <= x"10";
      when x"0814" => ROM_dataout_i <= x"ff";
      when x"0815" => ROM_dataout_i <= x"10";
      when x"0816" => ROM_dataout_i <= x"10";
      when x"0817" => ROM_dataout_i <= x"10";
      when x"0818" => ROM_dataout_i <= x"10";
      when x"0819" => ROM_dataout_i <= x"10";
      when x"081a" => ROM_dataout_i <= x"10";
      when x"081b" => ROM_dataout_i <= x"f0";
      when x"0823" => ROM_dataout_i <= x"1f";
      when x"0824" => ROM_dataout_i <= x"10";
      when x"0825" => ROM_dataout_i <= x"10";
      when x"0826" => ROM_dataout_i <= x"10";
      when x"0827" => ROM_dataout_i <= x"10";
      when x"0828" => ROM_dataout_i <= x"ff";
      when x"0829" => ROM_dataout_i <= x"ff";
      when x"082a" => ROM_dataout_i <= x"ff";
      when x"082b" => ROM_dataout_i <= x"ff";
      when x"082c" => ROM_dataout_i <= x"ff";
      when x"082d" => ROM_dataout_i <= x"ff";
      when x"082e" => ROM_dataout_i <= x"ff";
      when x"082f" => ROM_dataout_i <= x"ff";
      when x"0834" => ROM_dataout_i <= x"ff";
      when x"0835" => ROM_dataout_i <= x"ff";
      when x"0836" => ROM_dataout_i <= x"ff";
      when x"0837" => ROM_dataout_i <= x"ff";
      when x"0838" => ROM_dataout_i <= x"f0";
      when x"0839" => ROM_dataout_i <= x"f0";
      when x"083a" => ROM_dataout_i <= x"f0";
      when x"083b" => ROM_dataout_i <= x"f0";
      when x"083c" => ROM_dataout_i <= x"f0";
      when x"083d" => ROM_dataout_i <= x"f0";
      when x"083e" => ROM_dataout_i <= x"f0";
      when x"083f" => ROM_dataout_i <= x"f0";
      when x"0840" => ROM_dataout_i <= x"0f";
      when x"0841" => ROM_dataout_i <= x"0f";
      when x"0842" => ROM_dataout_i <= x"0f";
      when x"0843" => ROM_dataout_i <= x"0f";
      when x"0844" => ROM_dataout_i <= x"0f";
      when x"0845" => ROM_dataout_i <= x"0f";
      when x"0846" => ROM_dataout_i <= x"0f";
      when x"0847" => ROM_dataout_i <= x"0f";
      when x"0848" => ROM_dataout_i <= x"ff";
      when x"0849" => ROM_dataout_i <= x"ff";
      when x"084a" => ROM_dataout_i <= x"ff";
      when x"084b" => ROM_dataout_i <= x"ff";
      when x"0853" => ROM_dataout_i <= x"72";
      when x"0854" => ROM_dataout_i <= x"8c";
      when x"0855" => ROM_dataout_i <= x"88";
      when x"0856" => ROM_dataout_i <= x"3a";
      when x"0858" => ROM_dataout_i <= x"30";
      when x"0859" => ROM_dataout_i <= x"48";
      when x"085a" => ROM_dataout_i <= x"48";
      when x"085b" => ROM_dataout_i <= x"7c";
      when x"085c" => ROM_dataout_i <= x"42";
      when x"085d" => ROM_dataout_i <= x"42";
      when x"085e" => ROM_dataout_i <= x"dc";
      when x"0862" => ROM_dataout_i <= x"fe";
      when x"0863" => ROM_dataout_i <= x"42";
      when x"0864" => ROM_dataout_i <= x"40";
      when x"0865" => ROM_dataout_i <= x"40";
      when x"0866" => ROM_dataout_i <= x"e0";
      when x"086a" => ROM_dataout_i <= x"fe";
      when x"086b" => ROM_dataout_i <= x"44";
      when x"086c" => ROM_dataout_i <= x"44";
      when x"086d" => ROM_dataout_i <= x"44";
      when x"086e" => ROM_dataout_i <= x"ee";
      when x"0870" => ROM_dataout_i <= x"fe";
      when x"0871" => ROM_dataout_i <= x"42";
      when x"0872" => ROM_dataout_i <= x"20";
      when x"0873" => ROM_dataout_i <= x"10";
      when x"0874" => ROM_dataout_i <= x"20";
      when x"0875" => ROM_dataout_i <= x"42";
      when x"0876" => ROM_dataout_i <= x"fe";
      when x"087b" => ROM_dataout_i <= x"3e";
      when x"087c" => ROM_dataout_i <= x"44";
      when x"087d" => ROM_dataout_i <= x"44";
      when x"087e" => ROM_dataout_i <= x"38";
      when x"0882" => ROM_dataout_i <= x"cc";
      when x"0883" => ROM_dataout_i <= x"44";
      when x"0884" => ROM_dataout_i <= x"44";
      when x"0885" => ROM_dataout_i <= x"44";
      when x"0886" => ROM_dataout_i <= x"7a";
      when x"0887" => ROM_dataout_i <= x"40";
      when x"088a" => ROM_dataout_i <= x"7c";
      when x"088b" => ROM_dataout_i <= x"10";
      when x"088c" => ROM_dataout_i <= x"10";
      when x"088d" => ROM_dataout_i <= x"10";
      when x"088e" => ROM_dataout_i <= x"1c";
      when x"0891" => ROM_dataout_i <= x"10";
      when x"0892" => ROM_dataout_i <= x"7c";
      when x"0893" => ROM_dataout_i <= x"92";
      when x"0894" => ROM_dataout_i <= x"92";
      when x"0895" => ROM_dataout_i <= x"7c";
      when x"0896" => ROM_dataout_i <= x"10";
      when x"089a" => ROM_dataout_i <= x"7c";
      when x"089b" => ROM_dataout_i <= x"82";
      when x"089c" => ROM_dataout_i <= x"ba";
      when x"089d" => ROM_dataout_i <= x"82";
      when x"089e" => ROM_dataout_i <= x"7c";
      when x"08a3" => ROM_dataout_i <= x"7c";
      when x"08a4" => ROM_dataout_i <= x"82";
      when x"08a5" => ROM_dataout_i <= x"82";
      when x"08a6" => ROM_dataout_i <= x"6c";
      when x"08a7" => ROM_dataout_i <= x"28";
      when x"08a8" => ROM_dataout_i <= x"ee";
      when x"08ab" => ROM_dataout_i <= x"7c";
      when x"08ac" => ROM_dataout_i <= x"20";
      when x"08ad" => ROM_dataout_i <= x"38";
      when x"08ae" => ROM_dataout_i <= x"44";
      when x"08af" => ROM_dataout_i <= x"44";
      when x"08b0" => ROM_dataout_i <= x"38";
      when x"08b4" => ROM_dataout_i <= x"6c";
      when x"08b5" => ROM_dataout_i <= x"92";
      when x"08b6" => ROM_dataout_i <= x"92";
      when x"08b7" => ROM_dataout_i <= x"6c";
      when x"08bc" => ROM_dataout_i <= x"4c";
      when x"08bd" => ROM_dataout_i <= x"92";
      when x"08be" => ROM_dataout_i <= x"92";
      when x"08bf" => ROM_dataout_i <= x"7c";
      when x"08c0" => ROM_dataout_i <= x"10";
      when x"08c4" => ROM_dataout_i <= x"3c";
      when x"08c5" => ROM_dataout_i <= x"40";
      when x"08c6" => ROM_dataout_i <= x"30";
      when x"08c7" => ROM_dataout_i <= x"40";
      when x"08c8" => ROM_dataout_i <= x"3c";
      when x"08cc" => ROM_dataout_i <= x"3c";
      when x"08cd" => ROM_dataout_i <= x"42";
      when x"08ce" => ROM_dataout_i <= x"42";
      when x"08cf" => ROM_dataout_i <= x"42";
      when x"08d0" => ROM_dataout_i <= x"42";
      when x"08d3" => ROM_dataout_i <= x"fe";
      when x"08d5" => ROM_dataout_i <= x"fe";
      when x"08d7" => ROM_dataout_i <= x"fe";
      when x"08da" => ROM_dataout_i <= x"10";
      when x"08db" => ROM_dataout_i <= x"10";
      when x"08dc" => ROM_dataout_i <= x"fe";
      when x"08dd" => ROM_dataout_i <= x"10";
      when x"08de" => ROM_dataout_i <= x"10";
      when x"08df" => ROM_dataout_i <= x"fe";
      when x"08e2" => ROM_dataout_i <= x"40";
      when x"08e3" => ROM_dataout_i <= x"10";
      when x"08e4" => ROM_dataout_i <= x"04";
      when x"08e5" => ROM_dataout_i <= x"10";
      when x"08e6" => ROM_dataout_i <= x"40";
      when x"08e7" => ROM_dataout_i <= x"fe";
      when x"08ea" => ROM_dataout_i <= x"04";
      when x"08eb" => ROM_dataout_i <= x"10";
      when x"08ec" => ROM_dataout_i <= x"40";
      when x"08ed" => ROM_dataout_i <= x"10";
      when x"08ee" => ROM_dataout_i <= x"04";
      when x"08ef" => ROM_dataout_i <= x"fe";
      when x"08f2" => ROM_dataout_i <= x"0c";
      when x"08f3" => ROM_dataout_i <= x"10";
      when x"08f4" => ROM_dataout_i <= x"10";
      when x"08f5" => ROM_dataout_i <= x"10";
      when x"08f6" => ROM_dataout_i <= x"10";
      when x"08f7" => ROM_dataout_i <= x"10";
      when x"08f8" => ROM_dataout_i <= x"10";
      when x"08f9" => ROM_dataout_i <= x"10";
      when x"08fa" => ROM_dataout_i <= x"10";
      when x"08fb" => ROM_dataout_i <= x"10";
      when x"08fc" => ROM_dataout_i <= x"10";
      when x"08fd" => ROM_dataout_i <= x"10";
      when x"08fe" => ROM_dataout_i <= x"10";
      when x"08ff" => ROM_dataout_i <= x"10";
      when x"0900" => ROM_dataout_i <= x"10";
      when x"0901" => ROM_dataout_i <= x"60";
      when x"0904" => ROM_dataout_i <= x"10";
      when x"0906" => ROM_dataout_i <= x"fe";
      when x"0908" => ROM_dataout_i <= x"10";
      when x"090b" => ROM_dataout_i <= x"62";
      when x"090c" => ROM_dataout_i <= x"9c";
      when x"090e" => ROM_dataout_i <= x"62";
      when x"090f" => ROM_dataout_i <= x"9c";
      when x"0912" => ROM_dataout_i <= x"30";
      when x"0913" => ROM_dataout_i <= x"48";
      when x"0914" => ROM_dataout_i <= x"48";
      when x"0915" => ROM_dataout_i <= x"30";
      when x"091d" => ROM_dataout_i <= x"30";
      when x"091e" => ROM_dataout_i <= x"30";
      when x"0926" => ROM_dataout_i <= x"08";
      when x"092a" => ROM_dataout_i <= x"01";
      when x"092b" => ROM_dataout_i <= x"02";
      when x"092c" => ROM_dataout_i <= x"e2";
      when x"092d" => ROM_dataout_i <= x"24";
      when x"092e" => ROM_dataout_i <= x"14";
      when x"092f" => ROM_dataout_i <= x"18";
      when x"0930" => ROM_dataout_i <= x"08";
      when x"0934" => ROM_dataout_i <= x"58";
      when x"0935" => ROM_dataout_i <= x"24";
      when x"0936" => ROM_dataout_i <= x"24";
      when x"093a" => ROM_dataout_i <= x"30";
      when x"093b" => ROM_dataout_i <= x"48";
      when x"093c" => ROM_dataout_i <= x"10";
      when x"093d" => ROM_dataout_i <= x"20";
      when x"093e" => ROM_dataout_i <= x"78";
      when x"0944" => ROM_dataout_i <= x"ff";
      when x"0945" => ROM_dataout_i <= x"ff";
      when x"0946" => ROM_dataout_i <= x"ff";
      when x"0947" => ROM_dataout_i <= x"ff";
      when x"0953" => ROM_dataout_i <= x"f3";
      when x"0954" => ROM_dataout_i <= x"31";
      when x"0955" => ROM_dataout_i <= x"ff";
      when x"0956" => ROM_dataout_i <= x"ff";
      when x"0957" => ROM_dataout_i <= x"3e";
      when x"0958" => ROM_dataout_i <= x"e4";
      when x"0959" => ROM_dataout_i <= x"e0";
      when x"095a" => ROM_dataout_i <= x"47";
      when x"095b" => ROM_dataout_i <= x"3e";
      when x"095d" => ROM_dataout_i <= x"e0";
      when x"095e" => ROM_dataout_i <= x"43";
      when x"095f" => ROM_dataout_i <= x"e0";
      when x"0960" => ROM_dataout_i <= x"42";
      when x"0961" => ROM_dataout_i <= x"cd";
      when x"0962" => ROM_dataout_i <= x"9d";
      when x"0963" => ROM_dataout_i <= x"09";
      when x"0964" => ROM_dataout_i <= x"21";
      when x"0965" => ROM_dataout_i <= x"50";
      when x"0966" => ROM_dataout_i <= x"01";
      when x"0967" => ROM_dataout_i <= x"11";
      when x"0969" => ROM_dataout_i <= x"80";
      when x"096a" => ROM_dataout_i <= x"01";
      when x"096c" => ROM_dataout_i <= x"08";
      when x"096d" => ROM_dataout_i <= x"cd";
      when x"096e" => ROM_dataout_i <= x"7b";
      when x"0970" => ROM_dataout_i <= x"3e";
      when x"0971" => ROM_dataout_i <= x"95";
      when x"0972" => ROM_dataout_i <= x"e0";
      when x"0973" => ROM_dataout_i <= x"40";
      when x"0974" => ROM_dataout_i <= x"3e";
      when x"0975" => ROM_dataout_i <= x"20";
      when x"0976" => ROM_dataout_i <= x"21";
      when x"0978" => ROM_dataout_i <= x"98";
      when x"0979" => ROM_dataout_i <= x"01";
      when x"097b" => ROM_dataout_i <= x"04";
      when x"097c" => ROM_dataout_i <= x"cd";
      when x"097d" => ROM_dataout_i <= x"8b";
      when x"097f" => ROM_dataout_i <= x"21";
      when x"0980" => ROM_dataout_i <= x"90";
      when x"0981" => ROM_dataout_i <= x"09";
      when x"0982" => ROM_dataout_i <= x"11";
      when x"0983" => ROM_dataout_i <= x"e3";
      when x"0984" => ROM_dataout_i <= x"98";
      when x"0985" => ROM_dataout_i <= x"01";
      when x"0986" => ROM_dataout_i <= x"0d";
      when x"0988" => ROM_dataout_i <= x"cd";
      when x"0989" => ROM_dataout_i <= x"a1";
      when x"098b" => ROM_dataout_i <= x"76";
      when x"098e" => ROM_dataout_i <= x"18";
      when x"098f" => ROM_dataout_i <= x"fb";
      when x"0990" => ROM_dataout_i <= x"48";
      when x"0991" => ROM_dataout_i <= x"65";
      when x"0992" => ROM_dataout_i <= x"6c";
      when x"0993" => ROM_dataout_i <= x"6c";
      when x"0994" => ROM_dataout_i <= x"6f";
      when x"0995" => ROM_dataout_i <= x"20";
      when x"0996" => ROM_dataout_i <= x"57";
      when x"0997" => ROM_dataout_i <= x"6f";
      when x"0998" => ROM_dataout_i <= x"72";
      when x"0999" => ROM_dataout_i <= x"6c";
      when x"099a" => ROM_dataout_i <= x"64";
      when x"099b" => ROM_dataout_i <= x"20";
      when x"099c" => ROM_dataout_i <= x"21";
      when x"099d" => ROM_dataout_i <= x"f0";
      when x"099e" => ROM_dataout_i <= x"40";
      when x"099f" => ROM_dataout_i <= x"07";
      when x"09a0" => ROM_dataout_i <= x"d0";
      when x"09a1" => ROM_dataout_i <= x"f0";
      when x"09a2" => ROM_dataout_i <= x"44";
      when x"09a3" => ROM_dataout_i <= x"fe";
      when x"09a4" => ROM_dataout_i <= x"91";
      when x"09a5" => ROM_dataout_i <= x"20";
      when x"09a6" => ROM_dataout_i <= x"fa";
      when x"09a7" => ROM_dataout_i <= x"f0";
      when x"09a8" => ROM_dataout_i <= x"40";
      when x"09a9" => ROM_dataout_i <= x"cb";
      when x"09aa" => ROM_dataout_i <= x"bf";
      when x"09ab" => ROM_dataout_i <= x"e0";
      when x"09ac" => ROM_dataout_i <= x"40";
      when x"09ad" => ROM_dataout_i <= x"c9";
      when others => ROM_dataout_i <= x"00";
    end case;
  end process;


  --PREG: process(reset, clock)
  --begin
  --  if reset = '1' then 
  --    ROM_dataout <= x"00";
  --  elsif rising_edge(clock) then 
  --    ROM_dataout <= ROM_dataout_i;
  --  end if;
  --end process;
  ROM_dataout <= ROM_dataout_i;

  -------------------------------------------------------------------------------
  -- DEVICE UNDER TEST
  -------------------------------------------------------------------------------
  DUT: component processor port map(
    reset => reset,
    clock => clock,
    ROM_address => ROM_address,
    ROM_dataout => ROM_dataout);

  -------------------------------------------------------------------------------
  -- CLOCK
  -------------------------------------------------------------------------------
  PCLK: process
  begin
    clock <= '1';
    wait for clock_period/2;
    clock <= '0';
    wait for clock_period/2;
  end process;
  
end Behavioural;
